LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.my_inverse_pac.ALL;

ENTITY my_inverse IS
  PORT( clk                               :   IN    std_logic;
        reset_x                           :   IN    std_logic;
        clk_enable                        :   IN    std_logic;
        reset                             :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal1                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal2                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal3                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal4                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal5                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal6                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal7                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal8                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal9                   :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal10                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal11                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal12                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal13                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal14                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal15                  :   IN    std_logic_vector(7 DOWNTO 0);
        inBytes_signal16                  :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal1                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal2                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal3                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal4                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal5                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal6                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal7                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal8                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal9                       :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal10                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal11                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal12                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal13                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal14                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal15                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal16                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal17                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal18                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal19                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal20                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal21                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal22                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal23                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal24                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal25                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal26                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal27                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal28                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal29                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal30                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal31                      :   IN    std_logic_vector(7 DOWNTO 0);
        key_signal32                      :   IN    std_logic_vector(7 DOWNTO 0);
        ce_out                            :   OUT   std_logic;
        out_rsvd                          :   OUT   vector_of_std_logic_vector8(0 TO 15);
        valid                             :   OUT   std_logic_vector(7 DOWNTO 0);
        sit_out                           :   OUT   std_logic_vector(7 DOWNTO 0)
        );
END my_inverse;


ARCHITECTURE rtl OF my_inverse IS

  -- Signals
  SIGNAL enb                              : std_logic;
  SIGNAL reset_unsigned                   : unsigned(7 DOWNTO 0);
  SIGNAL Delay6_reg_rsvd                  : vector_of_unsigned8(0 TO 10);
  SIGNAL Delay6_reg_next                  : vector_of_unsigned8(0 TO 10);
  SIGNAL Delay6_out1                      : unsigned(7 DOWNTO 0);
  SIGNAL out0                             : std_logic;
  SIGNAL const_expression                 : unsigned(7 DOWNTO 0);
  SIGNAL sit                              : unsigned(7 DOWNTO 0);
  SIGNAL sit_1                            : unsigned(7 DOWNTO 0);
  SIGNAL ii                               : unsigned(7 DOWNTO 0);
  SIGNAL ii_1                             : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out          : std_logic;
  SIGNAL intdelay_ctrl_delay_out          : std_logic;
  SIGNAL intdelay_Initial_Val_out         : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_1               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_2               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_3               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_4               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_5               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_6               : unsigned(7 DOWNTO 0);
  SIGNAL ii_2                             : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_7               : unsigned(7 DOWNTO 0);
  SIGNAL sit_2                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_3                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_4                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_5                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_6                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_7                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_8                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_9                            : unsigned(7 DOWNTO 0);
  SIGNAL sit_10                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_11                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_1                           : std_logic;
  SIGNAL sit_12                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_2                           : std_logic;
  SIGNAL sit_13                           : unsigned(7 DOWNTO 0);
  SIGNAL ii_3                             : unsigned(7 DOWNTO 0);
  SIGNAL ii_4                             : unsigned(7 DOWNTO 0);
  SIGNAL i_i                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_3                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_4                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_5                           : std_logic;
  SIGNAL out0_6                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_7                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_8                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_9                           : std_logic;
  SIGNAL ii_5                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_10                          : std_logic;
  SIGNAL i_i_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_11                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_12                          : std_logic;
  SIGNAL out0_13                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_14                          : std_logic;
  SIGNAL out0_15                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_16                          : std_logic;
  SIGNAL out0_17                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_18                          : std_logic;
  SIGNAL out0_19                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_20                          : std_logic;
  SIGNAL out0_21                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_22                          : std_logic;
  SIGNAL out0_23                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_24                          : std_logic;
  SIGNAL i_i_2                            : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_out                     : unsigned(7 DOWNTO 0);
  SIGNAL ii_6                             : unsigned(7 DOWNTO 0);
  SIGNAL r_r                              : unsigned(7 DOWNTO 0);
  SIGNAL ii_7                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_25                          : unsigned(7 DOWNTO 0);
  SIGNAL ii_8                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_26                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_27                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_28                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_29                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_30                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_31                          : unsigned(7 DOWNTO 0);
  SIGNAL ii_9                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_32                          : std_logic;
  SIGNAL sit_14                           : unsigned(7 DOWNTO 0);
  SIGNAL sit_15                           : unsigned(7 DOWNTO 0);
  SIGNAL r_r_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_33                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_34                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_35                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_36                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_37                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_38                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_39                          : unsigned(7 DOWNTO 0);
  SIGNAL r_r_2                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_40                          : std_logic;
  SIGNAL sit_16                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_41                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_42                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_43                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_44                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_45                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_46                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_47                          : unsigned(7 DOWNTO 0);
  SIGNAL sit_out_1                        : unsigned(7 DOWNTO 0);
  SIGNAL sit_out_tmp                      : unsigned(7 DOWNTO 0);
  SIGNAL out0_48                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_49                          : unsigned(7 DOWNTO 0);
  SIGNAL j_j                              : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_8               : unsigned(7 DOWNTO 0);
  SIGNAL out0_50                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_9               : unsigned(7 DOWNTO 0);
  SIGNAL out0_51                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_10              : unsigned(7 DOWNTO 0);
  SIGNAL out0_52                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_11              : unsigned(7 DOWNTO 0);
  SIGNAL out0_53                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_12              : unsigned(7 DOWNTO 0);
  SIGNAL out0_54                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_13              : unsigned(15 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out_1        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_1        : std_logic;
  SIGNAL intdelay_Initial_Val_out_1       : vector_of_unsigned8(0 TO 255);
  SIGNAL sbox                             : vector_of_unsigned8(0 TO 255);
  SIGNAL intdelay_out_1                   : vector_of_unsigned8(0 TO 255);
  SIGNAL const_expression_14              : unsigned(15 DOWNTO 0);
  SIGNAL jj                               : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_15              : unsigned(7 DOWNTO 0);
  SIGNAL out0_55                          : unsigned(7 DOWNTO 0);
  SIGNAL iii                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_56                          : unsigned(7 DOWNTO 0);
  SIGNAL intdelay_ctrl_const_out_2        : std_logic;
  SIGNAL intdelay_ctrl_delay_out_2        : std_logic;
  SIGNAL intdelay_Initial_Val_out_2       : vector_of_unsigned8(0 TO 39);
  SIGNAL Rcon                             : vector_of_unsigned8(0 TO 39);
  SIGNAL intdelay_out_2                   : vector_of_unsigned8(0 TO 39);
  SIGNAL out0_57                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_16              : unsigned(7 DOWNTO 0);
  SIGNAL out0_58                          : unsigned(7 DOWNTO 0);
  SIGNAL iii_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_59                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_60                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_17              : unsigned(7 DOWNTO 0);
  SIGNAL out0_61                          : unsigned(7 DOWNTO 0);
  SIGNAL iii_2                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_62                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_63                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_18              : unsigned(7 DOWNTO 0);
  SIGNAL out0_64                          : unsigned(7 DOWNTO 0);
  SIGNAL iii_3                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_65                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_66                          : unsigned(7 DOWNTO 0);
  SIGNAL k2                               : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_67                          : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_1                             : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_2                             : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_68                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_69                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_70                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_71                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_72                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_73                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_74                          : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_3                             : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_4                             : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_5                             : vector_of_unsigned8(0 TO 3);
  SIGNAL k2_6                             : vector_of_unsigned8(0 TO 3);
  SIGNAL const_expression_19              : unsigned(7 DOWNTO 0);
  SIGNAL out0_75                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_20              : unsigned(7 DOWNTO 0);
  SIGNAL out0_76                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_21              : unsigned(7 DOWNTO 0);
  SIGNAL out0_77                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_22              : unsigned(7 DOWNTO 0);
  SIGNAL out0_78                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_23              : unsigned(7 DOWNTO 0);
  SIGNAL out0_79                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_24              : unsigned(7 DOWNTO 0);
  SIGNAL out0_80                          : unsigned(7 DOWNTO 0);
  SIGNAL const_expression_25              : unsigned(7 DOWNTO 0);
  SIGNAL out0_81                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal1_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal1                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal2_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal2                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal3_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal3                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal4_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal4                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal5_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal5                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal6_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal6                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal7_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal7                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal8_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal8                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal9_unsigned             : unsigned(7 DOWNTO 0);
  SIGNAL signal9                          : unsigned(7 DOWNTO 0);
  SIGNAL key_signal10_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal10                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal11_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal11                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal12_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal12                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal13_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal13                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal14_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal14                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal15_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal15                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal16_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal16                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal17_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal17                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal18_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal18                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal19_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal19                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal20_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal20                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal21_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal21                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal22_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal22                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal23_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal23                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal24_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal24                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal25_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal25                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal26_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal26                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal27_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal27                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal28_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal28                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal29_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal29                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal30_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal30                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal31_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal31                         : unsigned(7 DOWNTO 0);
  SIGNAL key_signal32_unsigned            : unsigned(7 DOWNTO 0);
  SIGNAL signal32                         : unsigned(7 DOWNTO 0);
  SIGNAL Delay5_out1_to_vector            : vector_of_unsigned8(0 TO 31);
  SIGNAL expandedKey                      : vector_of_unsigned8(0 TO 239);
  SIGNAL expandedKey_1                    : vector_of_unsigned8(0 TO 239);
  SIGNAL temp_key                         : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_3                       : unsigned(7 DOWNTO 0);
  SIGNAL expandedKey_2                    : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_82                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_83                          : unsigned(7 DOWNTO 0);
  SIGNAL temp_key_2                       : unsigned(7 DOWNTO 0);
  SIGNAL expandedKey_3                    : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_84                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_85                          : unsigned(7 DOWNTO 0);
  SIGNAL temp_key_1                       : unsigned(7 DOWNTO 0);
  SIGNAL expandedKey_4                    : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_86                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_87                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_88                          : vector_of_unsigned16(0 TO 3);
  SIGNAL out0_3_1                         : unsigned(15 DOWNTO 0);
  SIGNAL k1_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_2_1                         : unsigned(15 DOWNTO 0);
  SIGNAL k1_2                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_1_1                         : unsigned(15 DOWNTO 0);
  SIGNAL k1_1                             : unsigned(7 DOWNTO 0);
  SIGNAL temp_key_4                       : vector_of_unsigned8(0 TO 3);
  SIGNAL rotated_key                      : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_89                          : vector_of_unsigned16(0 TO 3);
  SIGNAL out0_0                           : unsigned(15 DOWNTO 0);
  SIGNAL k1_0                             : unsigned(7 DOWNTO 0);
  SIGNAL k1                               : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_5                       : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_90                          : vector_of_unsigned16(0 TO 3);
  SIGNAL out0_3_2                         : unsigned(15 DOWNTO 0);
  SIGNAL temp_key_3_1                     : unsigned(7 DOWNTO 0);
  SIGNAL out0_2_2                         : unsigned(15 DOWNTO 0);
  SIGNAL temp_key_2_1                     : unsigned(7 DOWNTO 0);
  SIGNAL out0_1_2                         : unsigned(15 DOWNTO 0);
  SIGNAL temp_key_1_1                     : unsigned(7 DOWNTO 0);
  SIGNAL out0_91                          : vector_of_unsigned16(0 TO 3);
  SIGNAL out0_0_1                         : unsigned(15 DOWNTO 0);
  SIGNAL temp_key_0                       : unsigned(7 DOWNTO 0);
  SIGNAL temp_key_6                       : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_92                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_93                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_94                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_95                          : unsigned(7 DOWNTO 0);
  SIGNAL temp_key_7                       : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_96                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_97                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_98                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_99                          : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_100                         : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_101                         : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_102                         : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_8                       : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_9                       : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_10                      : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_11                      : vector_of_unsigned8(0 TO 3);
  SIGNAL out0_103                         : vector_of_unsigned8(0 TO 3);
  SIGNAL temp_key_0_1                     : unsigned(7 DOWNTO 0);
  SIGNAL out0_104                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_105                         : unsigned(7 DOWNTO 0);
  SIGNAL expandedKey_5                    : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_106                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_107                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_108                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_109                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_110                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_111                         : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_112                         : vector_of_unsigned8(0 TO 239);
  SIGNAL expandedKey_6                    : vector_of_unsigned8(0 TO 239);
  SIGNAL out0_113                         : unsigned(7 DOWNTO 0);
  SIGNAL ss                               : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_114                         : vector_of_unsigned8(0 TO 15);
  SIGNAL ss_1                             : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_115                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_116                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_117                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_118                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_119                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_120                         : vector_of_unsigned8(0 TO 15);
  SIGNAL ss_2                             : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_121                         : unsigned(7 DOWNTO 0);
  SIGNAL gmul2                            : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3                            : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_1                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_1                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_2                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_2                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_3                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_3                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_4                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_4                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_5                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_5                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_6                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_6                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_7                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_7                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_8                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_8                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_9                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_9                          : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_10                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_10                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_11                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_11                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_12                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_12                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_13                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_13                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_14                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_14                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul3_15                         : vector_of_unsigned8(0 TO 255);
  SIGNAL gmul2_15                         : vector_of_unsigned8(0 TO 255);
  SIGNAL const_expression_26              : unsigned(15 DOWNTO 0);
  SIGNAL out0_122                         : vector_of_unsigned8(0 TO 15);
  SIGNAL inBytes_signal1_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal1_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal2_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal2_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal3_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal3_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal4_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal4_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal5_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal5_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal6_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal6_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal7_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal7_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal8_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal8_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal9_unsigned         : unsigned(7 DOWNTO 0);
  SIGNAL signal9_1                        : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal10_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal10_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal11_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal11_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal12_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal12_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal13_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal13_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal14_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal14_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal15_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal15_1                       : unsigned(7 DOWNTO 0);
  SIGNAL inBytes_signal16_unsigned        : unsigned(7 DOWNTO 0);
  SIGNAL signal16_1                       : unsigned(7 DOWNTO 0);
  SIGNAL Delay1_out1_to_vector            : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s                              : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_1                            : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_123                         : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_2                            : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_124                         : vector_of_unsigned16(0 TO 15);
  SIGNAL out0_11_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_11                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_6_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_6                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_1_3                         : unsigned(15 DOWNTO 0);
  SIGNAL s_1                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_12_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_12                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_7_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_7                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_2_3                         : unsigned(15 DOWNTO 0);
  SIGNAL s_2                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_13_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_13                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_8_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_8                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_3_3                         : unsigned(15 DOWNTO 0);
  SIGNAL s_3                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_14_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_14                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_9_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_9                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_4_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_4                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_15_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_15                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_10_1                        : unsigned(15 DOWNTO 0);
  SIGNAL s_10                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_5_1                         : unsigned(15 DOWNTO 0);
  SIGNAL s_5                              : unsigned(7 DOWNTO 0);
  SIGNAL out0_125                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_126                         : vector_of_unsigned16(0 TO 15);
  SIGNAL out0_0_2                         : unsigned(15 DOWNTO 0);
  SIGNAL s_0                              : unsigned(7 DOWNTO 0);
  SIGNAL s_s_3                            : vector_of_unsigned8(0 TO 15);
  SIGNAL s_15_1                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_127                         : unsigned(7 DOWNTO 0);
  SIGNAL s_12_1                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_128                         : unsigned(7 DOWNTO 0);
  SIGNAL s_13_1                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_129                         : unsigned(7 DOWNTO 0);
  SIGNAL s_14_1                           : unsigned(7 DOWNTO 0);
  SIGNAL b4                               : unsigned(7 DOWNTO 0);
  SIGNAL out0_130                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_131                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_132                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_133                         : unsigned(7 DOWNTO 0);
  SIGNAL b3                               : unsigned(7 DOWNTO 0);
  SIGNAL out0_134                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_135                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_136                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_137                         : unsigned(7 DOWNTO 0);
  SIGNAL b2                               : unsigned(7 DOWNTO 0);
  SIGNAL out0_138                         : unsigned(7 DOWNTO 0);
  SIGNAL s_s_4                            : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_139                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_140                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_141                         : unsigned(7 DOWNTO 0);
  SIGNAL b1                               : unsigned(7 DOWNTO 0);
  SIGNAL out0_142                         : unsigned(7 DOWNTO 0);
  SIGNAL s_11_1                           : unsigned(7 DOWNTO 0);
  SIGNAL out0_143                         : unsigned(7 DOWNTO 0);
  SIGNAL s_8_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_144                         : unsigned(7 DOWNTO 0);
  SIGNAL s_9_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_145                         : unsigned(7 DOWNTO 0);
  SIGNAL s_10_1                           : unsigned(7 DOWNTO 0);
  SIGNAL b4_1                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_146                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_147                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_148                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_149                         : unsigned(7 DOWNTO 0);
  SIGNAL b3_1                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_150                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_151                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_152                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_153                         : unsigned(7 DOWNTO 0);
  SIGNAL b2_1                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_154                         : unsigned(7 DOWNTO 0);
  SIGNAL s_s_5                            : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_155                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_156                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_157                         : unsigned(7 DOWNTO 0);
  SIGNAL b1_1                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_158                         : unsigned(7 DOWNTO 0);
  SIGNAL s_7_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_159                         : unsigned(7 DOWNTO 0);
  SIGNAL s_4_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_160                         : unsigned(7 DOWNTO 0);
  SIGNAL s_5_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_161                         : unsigned(7 DOWNTO 0);
  SIGNAL s_6_1                            : unsigned(7 DOWNTO 0);
  SIGNAL b4_2                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_162                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_163                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_164                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_165                         : unsigned(7 DOWNTO 0);
  SIGNAL b3_2                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_166                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_167                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_168                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_169                         : unsigned(7 DOWNTO 0);
  SIGNAL b2_2                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_170                         : unsigned(7 DOWNTO 0);
  SIGNAL s_s_6                            : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_171                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_172                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_173                         : unsigned(7 DOWNTO 0);
  SIGNAL b1_2                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_174                         : unsigned(7 DOWNTO 0);
  SIGNAL s_3_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_175                         : unsigned(7 DOWNTO 0);
  SIGNAL s_0_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_176                         : unsigned(7 DOWNTO 0);
  SIGNAL s_1_1                            : unsigned(7 DOWNTO 0);
  SIGNAL out0_177                         : unsigned(7 DOWNTO 0);
  SIGNAL s_2_1                            : unsigned(7 DOWNTO 0);
  SIGNAL b4_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_178                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_179                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_180                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_181                         : unsigned(7 DOWNTO 0);
  SIGNAL b3_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_182                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_183                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_184                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_185                         : unsigned(7 DOWNTO 0);
  SIGNAL b2_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_186                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_187                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_188                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_189                         : unsigned(7 DOWNTO 0);
  SIGNAL b1_3                             : unsigned(7 DOWNTO 0);
  SIGNAL out0_190                         : unsigned(7 DOWNTO 0);
  SIGNAL s_s_7                            : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_8                            : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_9                            : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_10                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_11                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_12                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_13                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_14                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_15                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_16                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_17                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_18                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_19                           : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_191                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_192                         : unsigned(7 DOWNTO 0);
  SIGNAL s_s_20                           : vector_of_unsigned8(0 TO 15);
  SIGNAL s_s_21                           : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_193                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_194                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_195                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_196                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_197                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_198                         : vector_of_unsigned8(0 TO 15);
  SIGNAL out0_199                         : vector_of_unsigned8(0 TO 15);
  SIGNAL Delay2_out1                      : vector_of_unsigned8(0 TO 15);
  SIGNAL valid_1                          : unsigned(7 DOWNTO 0);
  SIGNAL valid_2                          : unsigned(7 DOWNTO 0);
  SIGNAL valid_3                          : unsigned(7 DOWNTO 0);
  SIGNAL valid_4                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_200                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_5                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_201                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_6                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_202                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_7                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_203                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_8                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_204                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_9                          : unsigned(7 DOWNTO 0);
  SIGNAL out0_205                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_10                         : unsigned(7 DOWNTO 0);
  SIGNAL out0_206                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_11                         : unsigned(7 DOWNTO 0);
  SIGNAL valid_12                         : unsigned(7 DOWNTO 0);
  SIGNAL Delay3_out1                      : unsigned(7 DOWNTO 0);

BEGIN
  reset_unsigned <= unsigned(reset);

  enb <= clk_enable;

  Delay6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay6_reg_rsvd(0) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(1) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(2) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(3) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(4) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(5) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(6) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(7) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(8) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(9) <= to_unsigned(16#00#, 8);
        Delay6_reg_rsvd(10) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay6_reg_rsvd(0) <= Delay6_reg_next(0);
        Delay6_reg_rsvd(1) <= Delay6_reg_next(1);
        Delay6_reg_rsvd(2) <= Delay6_reg_next(2);
        Delay6_reg_rsvd(3) <= Delay6_reg_next(3);
        Delay6_reg_rsvd(4) <= Delay6_reg_next(4);
        Delay6_reg_rsvd(5) <= Delay6_reg_next(5);
        Delay6_reg_rsvd(6) <= Delay6_reg_next(6);
        Delay6_reg_rsvd(7) <= Delay6_reg_next(7);
        Delay6_reg_rsvd(8) <= Delay6_reg_next(8);
        Delay6_reg_rsvd(9) <= Delay6_reg_next(9);
        Delay6_reg_rsvd(10) <= Delay6_reg_next(10);
      END IF;
    END IF;
  END PROCESS Delay6_process;

  Delay6_out1 <= Delay6_reg_rsvd(10);
  Delay6_reg_next(0) <= reset_unsigned;
  Delay6_reg_next(1) <= Delay6_reg_rsvd(0);
  Delay6_reg_next(2) <= Delay6_reg_rsvd(1);
  Delay6_reg_next(3) <= Delay6_reg_rsvd(2);
  Delay6_reg_next(4) <= Delay6_reg_rsvd(3);
  Delay6_reg_next(5) <= Delay6_reg_rsvd(4);
  Delay6_reg_next(6) <= Delay6_reg_rsvd(5);
  Delay6_reg_next(7) <= Delay6_reg_rsvd(6);
  Delay6_reg_next(8) <= Delay6_reg_rsvd(7);
  Delay6_reg_next(9) <= Delay6_reg_rsvd(8);
  Delay6_reg_next(10) <= Delay6_reg_rsvd(9);

  
  out0 <= '1' WHEN Delay6_out1 = to_unsigned(16#01#, 8) ELSE
      '0';

  const_expression <= to_unsigned(16#01#, 8);

  sit <= to_unsigned(16#04#, 8);

  sit_1 <= to_unsigned(16#0E#, 8);

  ii <= to_unsigned(16#00#, 8);

  ii_1 <= to_unsigned(16#00#, 8);

  intdelay_ctrl_const_out <= '1';

  intdelay_ctrl_delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out <= intdelay_ctrl_const_out;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay2_process;


  intdelay_Initial_Val_out <= to_unsigned(16#08#, 8);

  const_expression_1 <= to_unsigned(16#01#, 8);

  const_expression_2 <= to_unsigned(16#01#, 8);

  const_expression_3 <= to_unsigned(16#07#, 8);

  const_expression_4 <= to_unsigned(16#01#, 8);

  const_expression_5 <= to_unsigned(16#07#, 8);

  const_expression_6 <= to_unsigned(16#01#, 8);

  ii_2 <= to_unsigned(16#01#, 8);

  const_expression_7 <= to_unsigned(16#01#, 8);

  sit_2 <= to_unsigned(16#0A#, 8);

  sit_3 <= to_unsigned(16#07#, 8);

  sit_4 <= to_unsigned(16#07#, 8);

  sit_5 <= to_unsigned(16#06#, 8);

  sit_6 <= to_unsigned(16#05#, 8);

  sit_7 <= to_unsigned(16#04#, 8);

  sit_8 <= to_unsigned(16#02#, 8);

  sit_9 <= to_unsigned(16#03#, 8);

  sit_10 <= to_unsigned(16#02#, 8);

  sit_11 <= to_unsigned(16#01#, 8);

  
  sit_12 <= sit_8 WHEN out0_1 = '0' ELSE
      sit_9;

  
  sit_13 <= sit_4 WHEN out0_2 = '0' ELSE
      sit_5;

  ii_4 <= ii_3 + const_expression_6;

  out0_3 <= i_i - const_expression_4;

  out0_4 <= out0_3 AND const_expression_5;

  
  out0_5 <= '1' WHEN out0_4 = to_unsigned(16#04#, 8) ELSE
      '0';

  
  out0_6 <= ii_3 WHEN out0_5 = '0' ELSE
      ii_3;

  out0_7 <= i_i - const_expression_2;

  out0_8 <= out0_7 AND const_expression_3;

  
  out0_9 <= '1' WHEN out0_8 = to_unsigned(16#00#, 8) ELSE
      '0';

  
  ii_5 <= out0_6 WHEN out0_9 = '0' ELSE
      ii_4;

  
  out0_11 <= i_i_1 WHEN out0_10 = '0' ELSE
      i_i_1;

  
  out0_13 <= out0_11 WHEN out0_12 = '0' ELSE
      i_i_1;

  
  out0_15 <= out0_13 WHEN out0_14 = '0' ELSE
      i_i_1;

  
  out0_17 <= out0_15 WHEN out0_16 = '0' ELSE
      i_i_1;

  
  out0_19 <= out0_17 WHEN out0_18 = '0' ELSE
      i_i_1;

  
  out0_21 <= out0_19 WHEN out0_20 = '0' ELSE
      i_i_1;

  
  out0_23 <= out0_21 WHEN out0_22 = '0' ELSE
      i_i;

  
  i_i_2 <= out0_23 WHEN out0_24 = '0' ELSE
      i_i_1;

  intdelay6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out <= i_i_2;
      END IF;
    END IF;
  END PROCESS intdelay6_process;


  
  i_i_1 <= intdelay_Initial_Val_out WHEN intdelay_ctrl_delay_out = '0' ELSE
      intdelay_out;

  i_i <= i_i_1 + const_expression_1;

  
  out0_1 <= '1' WHEN i_i = to_unsigned(16#3C#, 8) ELSE
      '0';

  
  ii_6 <= ii_5 WHEN out0_1 = '0' ELSE
      ii_2;

  
  out0_2 <= '1' WHEN r_r <= to_unsigned(16#0D#, 8) ELSE
      '0';

  
  ii_7 <= ii_1 WHEN out0_2 = '0' ELSE
      ii_3;

  
  out0_25 <= ii_3 WHEN out0_10 = '0' ELSE
      ii_3;

  
  out0_26 <= out0_25 WHEN out0_12 = '0' ELSE
      ii_8;

  
  out0_27 <= out0_26 WHEN out0_14 = '0' ELSE
      ii;

  
  out0_28 <= out0_27 WHEN out0_16 = '0' ELSE
      ii_7;

  
  out0_29 <= out0_28 WHEN out0_18 = '0' ELSE
      ii_3;

  
  out0_30 <= out0_29 WHEN out0_20 = '0' ELSE
      ii_3;

  
  out0_31 <= out0_30 WHEN out0_22 = '0' ELSE
      ii_6;

  
  ii_9 <= out0_31 WHEN out0_24 = '0' ELSE
      ii_3;

  intdelay7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        ii_3 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        ii_3 <= ii_9;
      END IF;
    END IF;
  END PROCESS intdelay7_process;


  ii_8 <= ii_3 + const_expression_7;

  
  out0_32 <= '1' WHEN ii_8 = to_unsigned(16#10#, 8) ELSE
      '0';

  
  sit_15 <= sit_14 WHEN out0_32 = '0' ELSE
      sit_2;

  r_r_1 <= r_r + const_expression;

  
  out0_33 <= r_r WHEN out0_10 = '0' ELSE
      r_r;

  
  out0_34 <= out0_33 WHEN out0_12 = '0' ELSE
      r_r;

  
  out0_35 <= out0_34 WHEN out0_14 = '0' ELSE
      r_r;

  
  out0_36 <= out0_35 WHEN out0_16 = '0' ELSE
      r_r;

  
  out0_37 <= out0_36 WHEN out0_18 = '0' ELSE
      r_r_1;

  
  out0_38 <= out0_37 WHEN out0_20 = '0' ELSE
      r_r;

  
  out0_39 <= out0_38 WHEN out0_22 = '0' ELSE
      r_r;

  
  r_r_2 <= out0_39 WHEN out0_24 = '0' ELSE
      r_r;

  intdelay8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        r_r <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        r_r <= r_r_2;
      END IF;
    END IF;
  END PROCESS intdelay8_process;


  
  out0_40 <= '1' WHEN r_r = to_unsigned(16#0E#, 8) ELSE
      '0';

  
  sit_16 <= sit WHEN out0_40 = '0' ELSE
      sit_1;

  
  out0_10 <= '1' WHEN sit_14 = to_unsigned(16#0A#, 8) ELSE
      '0';

  
  out0_41 <= sit_14 WHEN out0_10 = '0' ELSE
      sit_16;

  
  out0_12 <= '1' WHEN sit_14 = to_unsigned(16#07#, 8) ELSE
      '0';

  
  out0_42 <= out0_41 WHEN out0_12 = '0' ELSE
      sit_15;

  
  out0_14 <= '1' WHEN sit_14 = to_unsigned(16#06#, 8) ELSE
      '0';

  
  out0_43 <= out0_42 WHEN out0_14 = '0' ELSE
      sit_3;

  
  out0_16 <= '1' WHEN sit_14 = to_unsigned(16#05#, 8) ELSE
      '0';

  
  out0_44 <= out0_43 WHEN out0_16 = '0' ELSE
      sit_13;

  
  out0_18 <= '1' WHEN sit_14 = to_unsigned(16#04#, 8) ELSE
      '0';

  
  out0_45 <= out0_44 WHEN out0_18 = '0' ELSE
      sit_6;

  
  out0_20 <= '1' WHEN sit_14 = to_unsigned(16#03#, 8) ELSE
      '0';

  
  out0_46 <= out0_45 WHEN out0_20 = '0' ELSE
      sit_7;

  
  out0_22 <= '1' WHEN sit_14 = to_unsigned(16#02#, 8) ELSE
      '0';

  
  out0_47 <= out0_46 WHEN out0_22 = '0' ELSE
      sit_12;

  
  sit_out_1 <= out0_47 WHEN out0_24 = '0' ELSE
      sit_10;

  reduced_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        sit_out_tmp <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        sit_out_tmp <= sit_out_1;
      END IF;
    END IF;
  END PROCESS reduced_process;


  -- %
  
  sit_14 <= sit_out_tmp WHEN out0 = '0' ELSE
      sit_11;

  
  out0_24 <= '1' WHEN sit_14 = to_unsigned(16#01#, 8) ELSE
      '0';

  out0_48 <= r_r sll 4;

  out0_49 <= out0_48 + ii_8;

  j_j <= i_i sll 2;

  const_expression_8 <= to_unsigned(16#23#, 8);

  out0_50 <= j_j - const_expression_8;

  const_expression_9 <= to_unsigned(16#07#, 8);

  out0_51 <= j_j - const_expression_9;

  const_expression_10 <= to_unsigned(16#06#, 8);

  out0_52 <= j_j - const_expression_10;

  const_expression_11 <= to_unsigned(16#05#, 8);

  out0_53 <= j_j - const_expression_11;

  const_expression_12 <= to_unsigned(16#04#, 8);

  out0_54 <= j_j - const_expression_12;

  const_expression_13 <= to_unsigned(16#0001#, 16);

  intdelay_ctrl_const_out_1 <= '1';

  intdelay_ctrl_delay_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_1 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_1 <= intdelay_ctrl_const_out_1;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay_process;


  intdelay_Initial_Val_out_1(0) <= to_unsigned(16#63#, 8);
  intdelay_Initial_Val_out_1(1) <= to_unsigned(16#7C#, 8);
  intdelay_Initial_Val_out_1(2) <= to_unsigned(16#77#, 8);
  intdelay_Initial_Val_out_1(3) <= to_unsigned(16#7B#, 8);
  intdelay_Initial_Val_out_1(4) <= to_unsigned(16#F2#, 8);
  intdelay_Initial_Val_out_1(5) <= to_unsigned(16#6B#, 8);
  intdelay_Initial_Val_out_1(6) <= to_unsigned(16#6F#, 8);
  intdelay_Initial_Val_out_1(7) <= to_unsigned(16#C5#, 8);
  intdelay_Initial_Val_out_1(8) <= to_unsigned(16#30#, 8);
  intdelay_Initial_Val_out_1(9) <= to_unsigned(16#01#, 8);
  intdelay_Initial_Val_out_1(10) <= to_unsigned(16#67#, 8);
  intdelay_Initial_Val_out_1(11) <= to_unsigned(16#2B#, 8);
  intdelay_Initial_Val_out_1(12) <= to_unsigned(16#FE#, 8);
  intdelay_Initial_Val_out_1(13) <= to_unsigned(16#D7#, 8);
  intdelay_Initial_Val_out_1(14) <= to_unsigned(16#AB#, 8);
  intdelay_Initial_Val_out_1(15) <= to_unsigned(16#76#, 8);
  intdelay_Initial_Val_out_1(16) <= to_unsigned(16#CA#, 8);
  intdelay_Initial_Val_out_1(17) <= to_unsigned(16#82#, 8);
  intdelay_Initial_Val_out_1(18) <= to_unsigned(16#C9#, 8);
  intdelay_Initial_Val_out_1(19) <= to_unsigned(16#7D#, 8);
  intdelay_Initial_Val_out_1(20) <= to_unsigned(16#FA#, 8);
  intdelay_Initial_Val_out_1(21) <= to_unsigned(16#59#, 8);
  intdelay_Initial_Val_out_1(22) <= to_unsigned(16#47#, 8);
  intdelay_Initial_Val_out_1(23) <= to_unsigned(16#F0#, 8);
  intdelay_Initial_Val_out_1(24) <= to_unsigned(16#AD#, 8);
  intdelay_Initial_Val_out_1(25) <= to_unsigned(16#D4#, 8);
  intdelay_Initial_Val_out_1(26) <= to_unsigned(16#A2#, 8);
  intdelay_Initial_Val_out_1(27) <= to_unsigned(16#AF#, 8);
  intdelay_Initial_Val_out_1(28) <= to_unsigned(16#9C#, 8);
  intdelay_Initial_Val_out_1(29) <= to_unsigned(16#A4#, 8);
  intdelay_Initial_Val_out_1(30) <= to_unsigned(16#72#, 8);
  intdelay_Initial_Val_out_1(31) <= to_unsigned(16#C0#, 8);
  intdelay_Initial_Val_out_1(32) <= to_unsigned(16#B7#, 8);
  intdelay_Initial_Val_out_1(33) <= to_unsigned(16#FD#, 8);
  intdelay_Initial_Val_out_1(34) <= to_unsigned(16#93#, 8);
  intdelay_Initial_Val_out_1(35) <= to_unsigned(16#26#, 8);
  intdelay_Initial_Val_out_1(36) <= to_unsigned(16#36#, 8);
  intdelay_Initial_Val_out_1(37) <= to_unsigned(16#3F#, 8);
  intdelay_Initial_Val_out_1(38) <= to_unsigned(16#F7#, 8);
  intdelay_Initial_Val_out_1(39) <= to_unsigned(16#CC#, 8);
  intdelay_Initial_Val_out_1(40) <= to_unsigned(16#34#, 8);
  intdelay_Initial_Val_out_1(41) <= to_unsigned(16#A5#, 8);
  intdelay_Initial_Val_out_1(42) <= to_unsigned(16#E5#, 8);
  intdelay_Initial_Val_out_1(43) <= to_unsigned(16#F1#, 8);
  intdelay_Initial_Val_out_1(44) <= to_unsigned(16#71#, 8);
  intdelay_Initial_Val_out_1(45) <= to_unsigned(16#D8#, 8);
  intdelay_Initial_Val_out_1(46) <= to_unsigned(16#31#, 8);
  intdelay_Initial_Val_out_1(47) <= to_unsigned(16#15#, 8);
  intdelay_Initial_Val_out_1(48) <= to_unsigned(16#04#, 8);
  intdelay_Initial_Val_out_1(49) <= to_unsigned(16#C7#, 8);
  intdelay_Initial_Val_out_1(50) <= to_unsigned(16#23#, 8);
  intdelay_Initial_Val_out_1(51) <= to_unsigned(16#C3#, 8);
  intdelay_Initial_Val_out_1(52) <= to_unsigned(16#18#, 8);
  intdelay_Initial_Val_out_1(53) <= to_unsigned(16#96#, 8);
  intdelay_Initial_Val_out_1(54) <= to_unsigned(16#05#, 8);
  intdelay_Initial_Val_out_1(55) <= to_unsigned(16#9A#, 8);
  intdelay_Initial_Val_out_1(56) <= to_unsigned(16#07#, 8);
  intdelay_Initial_Val_out_1(57) <= to_unsigned(16#12#, 8);
  intdelay_Initial_Val_out_1(58) <= to_unsigned(16#80#, 8);
  intdelay_Initial_Val_out_1(59) <= to_unsigned(16#E2#, 8);
  intdelay_Initial_Val_out_1(60) <= to_unsigned(16#EB#, 8);
  intdelay_Initial_Val_out_1(61) <= to_unsigned(16#27#, 8);
  intdelay_Initial_Val_out_1(62) <= to_unsigned(16#B2#, 8);
  intdelay_Initial_Val_out_1(63) <= to_unsigned(16#75#, 8);
  intdelay_Initial_Val_out_1(64) <= to_unsigned(16#09#, 8);
  intdelay_Initial_Val_out_1(65) <= to_unsigned(16#83#, 8);
  intdelay_Initial_Val_out_1(66) <= to_unsigned(16#2C#, 8);
  intdelay_Initial_Val_out_1(67) <= to_unsigned(16#1A#, 8);
  intdelay_Initial_Val_out_1(68) <= to_unsigned(16#1B#, 8);
  intdelay_Initial_Val_out_1(69) <= to_unsigned(16#6E#, 8);
  intdelay_Initial_Val_out_1(70) <= to_unsigned(16#5A#, 8);
  intdelay_Initial_Val_out_1(71) <= to_unsigned(16#A0#, 8);
  intdelay_Initial_Val_out_1(72) <= to_unsigned(16#52#, 8);
  intdelay_Initial_Val_out_1(73) <= to_unsigned(16#3B#, 8);
  intdelay_Initial_Val_out_1(74) <= to_unsigned(16#D6#, 8);
  intdelay_Initial_Val_out_1(75) <= to_unsigned(16#B3#, 8);
  intdelay_Initial_Val_out_1(76) <= to_unsigned(16#29#, 8);
  intdelay_Initial_Val_out_1(77) <= to_unsigned(16#E3#, 8);
  intdelay_Initial_Val_out_1(78) <= to_unsigned(16#2F#, 8);
  intdelay_Initial_Val_out_1(79) <= to_unsigned(16#84#, 8);
  intdelay_Initial_Val_out_1(80) <= to_unsigned(16#53#, 8);
  intdelay_Initial_Val_out_1(81) <= to_unsigned(16#D1#, 8);
  intdelay_Initial_Val_out_1(82) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_1(83) <= to_unsigned(16#ED#, 8);
  intdelay_Initial_Val_out_1(84) <= to_unsigned(16#20#, 8);
  intdelay_Initial_Val_out_1(85) <= to_unsigned(16#FC#, 8);
  intdelay_Initial_Val_out_1(86) <= to_unsigned(16#B1#, 8);
  intdelay_Initial_Val_out_1(87) <= to_unsigned(16#5B#, 8);
  intdelay_Initial_Val_out_1(88) <= to_unsigned(16#6A#, 8);
  intdelay_Initial_Val_out_1(89) <= to_unsigned(16#CB#, 8);
  intdelay_Initial_Val_out_1(90) <= to_unsigned(16#BE#, 8);
  intdelay_Initial_Val_out_1(91) <= to_unsigned(16#39#, 8);
  intdelay_Initial_Val_out_1(92) <= to_unsigned(16#4A#, 8);
  intdelay_Initial_Val_out_1(93) <= to_unsigned(16#4C#, 8);
  intdelay_Initial_Val_out_1(94) <= to_unsigned(16#58#, 8);
  intdelay_Initial_Val_out_1(95) <= to_unsigned(16#CF#, 8);
  intdelay_Initial_Val_out_1(96) <= to_unsigned(16#D0#, 8);
  intdelay_Initial_Val_out_1(97) <= to_unsigned(16#EF#, 8);
  intdelay_Initial_Val_out_1(98) <= to_unsigned(16#AA#, 8);
  intdelay_Initial_Val_out_1(99) <= to_unsigned(16#FB#, 8);
  intdelay_Initial_Val_out_1(100) <= to_unsigned(16#43#, 8);
  intdelay_Initial_Val_out_1(101) <= to_unsigned(16#4D#, 8);
  intdelay_Initial_Val_out_1(102) <= to_unsigned(16#33#, 8);
  intdelay_Initial_Val_out_1(103) <= to_unsigned(16#85#, 8);
  intdelay_Initial_Val_out_1(104) <= to_unsigned(16#45#, 8);
  intdelay_Initial_Val_out_1(105) <= to_unsigned(16#F9#, 8);
  intdelay_Initial_Val_out_1(106) <= to_unsigned(16#02#, 8);
  intdelay_Initial_Val_out_1(107) <= to_unsigned(16#7F#, 8);
  intdelay_Initial_Val_out_1(108) <= to_unsigned(16#50#, 8);
  intdelay_Initial_Val_out_1(109) <= to_unsigned(16#3C#, 8);
  intdelay_Initial_Val_out_1(110) <= to_unsigned(16#9F#, 8);
  intdelay_Initial_Val_out_1(111) <= to_unsigned(16#A8#, 8);
  intdelay_Initial_Val_out_1(112) <= to_unsigned(16#51#, 8);
  intdelay_Initial_Val_out_1(113) <= to_unsigned(16#A3#, 8);
  intdelay_Initial_Val_out_1(114) <= to_unsigned(16#40#, 8);
  intdelay_Initial_Val_out_1(115) <= to_unsigned(16#8F#, 8);
  intdelay_Initial_Val_out_1(116) <= to_unsigned(16#92#, 8);
  intdelay_Initial_Val_out_1(117) <= to_unsigned(16#9D#, 8);
  intdelay_Initial_Val_out_1(118) <= to_unsigned(16#38#, 8);
  intdelay_Initial_Val_out_1(119) <= to_unsigned(16#F5#, 8);
  intdelay_Initial_Val_out_1(120) <= to_unsigned(16#BC#, 8);
  intdelay_Initial_Val_out_1(121) <= to_unsigned(16#B6#, 8);
  intdelay_Initial_Val_out_1(122) <= to_unsigned(16#DA#, 8);
  intdelay_Initial_Val_out_1(123) <= to_unsigned(16#21#, 8);
  intdelay_Initial_Val_out_1(124) <= to_unsigned(16#10#, 8);
  intdelay_Initial_Val_out_1(125) <= to_unsigned(16#FF#, 8);
  intdelay_Initial_Val_out_1(126) <= to_unsigned(16#F3#, 8);
  intdelay_Initial_Val_out_1(127) <= to_unsigned(16#D2#, 8);
  intdelay_Initial_Val_out_1(128) <= to_unsigned(16#CD#, 8);
  intdelay_Initial_Val_out_1(129) <= to_unsigned(16#0C#, 8);
  intdelay_Initial_Val_out_1(130) <= to_unsigned(16#13#, 8);
  intdelay_Initial_Val_out_1(131) <= to_unsigned(16#EC#, 8);
  intdelay_Initial_Val_out_1(132) <= to_unsigned(16#5F#, 8);
  intdelay_Initial_Val_out_1(133) <= to_unsigned(16#97#, 8);
  intdelay_Initial_Val_out_1(134) <= to_unsigned(16#44#, 8);
  intdelay_Initial_Val_out_1(135) <= to_unsigned(16#17#, 8);
  intdelay_Initial_Val_out_1(136) <= to_unsigned(16#C4#, 8);
  intdelay_Initial_Val_out_1(137) <= to_unsigned(16#A7#, 8);
  intdelay_Initial_Val_out_1(138) <= to_unsigned(16#7E#, 8);
  intdelay_Initial_Val_out_1(139) <= to_unsigned(16#3D#, 8);
  intdelay_Initial_Val_out_1(140) <= to_unsigned(16#64#, 8);
  intdelay_Initial_Val_out_1(141) <= to_unsigned(16#5D#, 8);
  intdelay_Initial_Val_out_1(142) <= to_unsigned(16#19#, 8);
  intdelay_Initial_Val_out_1(143) <= to_unsigned(16#73#, 8);
  intdelay_Initial_Val_out_1(144) <= to_unsigned(16#60#, 8);
  intdelay_Initial_Val_out_1(145) <= to_unsigned(16#81#, 8);
  intdelay_Initial_Val_out_1(146) <= to_unsigned(16#4F#, 8);
  intdelay_Initial_Val_out_1(147) <= to_unsigned(16#DC#, 8);
  intdelay_Initial_Val_out_1(148) <= to_unsigned(16#22#, 8);
  intdelay_Initial_Val_out_1(149) <= to_unsigned(16#2A#, 8);
  intdelay_Initial_Val_out_1(150) <= to_unsigned(16#90#, 8);
  intdelay_Initial_Val_out_1(151) <= to_unsigned(16#88#, 8);
  intdelay_Initial_Val_out_1(152) <= to_unsigned(16#46#, 8);
  intdelay_Initial_Val_out_1(153) <= to_unsigned(16#EE#, 8);
  intdelay_Initial_Val_out_1(154) <= to_unsigned(16#B8#, 8);
  intdelay_Initial_Val_out_1(155) <= to_unsigned(16#14#, 8);
  intdelay_Initial_Val_out_1(156) <= to_unsigned(16#DE#, 8);
  intdelay_Initial_Val_out_1(157) <= to_unsigned(16#5E#, 8);
  intdelay_Initial_Val_out_1(158) <= to_unsigned(16#0B#, 8);
  intdelay_Initial_Val_out_1(159) <= to_unsigned(16#DB#, 8);
  intdelay_Initial_Val_out_1(160) <= to_unsigned(16#E0#, 8);
  intdelay_Initial_Val_out_1(161) <= to_unsigned(16#32#, 8);
  intdelay_Initial_Val_out_1(162) <= to_unsigned(16#3A#, 8);
  intdelay_Initial_Val_out_1(163) <= to_unsigned(16#0A#, 8);
  intdelay_Initial_Val_out_1(164) <= to_unsigned(16#49#, 8);
  intdelay_Initial_Val_out_1(165) <= to_unsigned(16#06#, 8);
  intdelay_Initial_Val_out_1(166) <= to_unsigned(16#24#, 8);
  intdelay_Initial_Val_out_1(167) <= to_unsigned(16#5C#, 8);
  intdelay_Initial_Val_out_1(168) <= to_unsigned(16#C2#, 8);
  intdelay_Initial_Val_out_1(169) <= to_unsigned(16#D3#, 8);
  intdelay_Initial_Val_out_1(170) <= to_unsigned(16#AC#, 8);
  intdelay_Initial_Val_out_1(171) <= to_unsigned(16#62#, 8);
  intdelay_Initial_Val_out_1(172) <= to_unsigned(16#91#, 8);
  intdelay_Initial_Val_out_1(173) <= to_unsigned(16#95#, 8);
  intdelay_Initial_Val_out_1(174) <= to_unsigned(16#E4#, 8);
  intdelay_Initial_Val_out_1(175) <= to_unsigned(16#79#, 8);
  intdelay_Initial_Val_out_1(176) <= to_unsigned(16#E7#, 8);
  intdelay_Initial_Val_out_1(177) <= to_unsigned(16#C8#, 8);
  intdelay_Initial_Val_out_1(178) <= to_unsigned(16#37#, 8);
  intdelay_Initial_Val_out_1(179) <= to_unsigned(16#6D#, 8);
  intdelay_Initial_Val_out_1(180) <= to_unsigned(16#8D#, 8);
  intdelay_Initial_Val_out_1(181) <= to_unsigned(16#D5#, 8);
  intdelay_Initial_Val_out_1(182) <= to_unsigned(16#4E#, 8);
  intdelay_Initial_Val_out_1(183) <= to_unsigned(16#A9#, 8);
  intdelay_Initial_Val_out_1(184) <= to_unsigned(16#6C#, 8);
  intdelay_Initial_Val_out_1(185) <= to_unsigned(16#56#, 8);
  intdelay_Initial_Val_out_1(186) <= to_unsigned(16#F4#, 8);
  intdelay_Initial_Val_out_1(187) <= to_unsigned(16#EA#, 8);
  intdelay_Initial_Val_out_1(188) <= to_unsigned(16#65#, 8);
  intdelay_Initial_Val_out_1(189) <= to_unsigned(16#7A#, 8);
  intdelay_Initial_Val_out_1(190) <= to_unsigned(16#AE#, 8);
  intdelay_Initial_Val_out_1(191) <= to_unsigned(16#08#, 8);
  intdelay_Initial_Val_out_1(192) <= to_unsigned(16#BA#, 8);
  intdelay_Initial_Val_out_1(193) <= to_unsigned(16#78#, 8);
  intdelay_Initial_Val_out_1(194) <= to_unsigned(16#25#, 8);
  intdelay_Initial_Val_out_1(195) <= to_unsigned(16#2E#, 8);
  intdelay_Initial_Val_out_1(196) <= to_unsigned(16#1C#, 8);
  intdelay_Initial_Val_out_1(197) <= to_unsigned(16#A6#, 8);
  intdelay_Initial_Val_out_1(198) <= to_unsigned(16#B4#, 8);
  intdelay_Initial_Val_out_1(199) <= to_unsigned(16#C6#, 8);
  intdelay_Initial_Val_out_1(200) <= to_unsigned(16#E8#, 8);
  intdelay_Initial_Val_out_1(201) <= to_unsigned(16#DD#, 8);
  intdelay_Initial_Val_out_1(202) <= to_unsigned(16#74#, 8);
  intdelay_Initial_Val_out_1(203) <= to_unsigned(16#1F#, 8);
  intdelay_Initial_Val_out_1(204) <= to_unsigned(16#4B#, 8);
  intdelay_Initial_Val_out_1(205) <= to_unsigned(16#BD#, 8);
  intdelay_Initial_Val_out_1(206) <= to_unsigned(16#8B#, 8);
  intdelay_Initial_Val_out_1(207) <= to_unsigned(16#8A#, 8);
  intdelay_Initial_Val_out_1(208) <= to_unsigned(16#70#, 8);
  intdelay_Initial_Val_out_1(209) <= to_unsigned(16#3E#, 8);
  intdelay_Initial_Val_out_1(210) <= to_unsigned(16#B5#, 8);
  intdelay_Initial_Val_out_1(211) <= to_unsigned(16#66#, 8);
  intdelay_Initial_Val_out_1(212) <= to_unsigned(16#48#, 8);
  intdelay_Initial_Val_out_1(213) <= to_unsigned(16#03#, 8);
  intdelay_Initial_Val_out_1(214) <= to_unsigned(16#F6#, 8);
  intdelay_Initial_Val_out_1(215) <= to_unsigned(16#0E#, 8);
  intdelay_Initial_Val_out_1(216) <= to_unsigned(16#61#, 8);
  intdelay_Initial_Val_out_1(217) <= to_unsigned(16#35#, 8);
  intdelay_Initial_Val_out_1(218) <= to_unsigned(16#57#, 8);
  intdelay_Initial_Val_out_1(219) <= to_unsigned(16#B9#, 8);
  intdelay_Initial_Val_out_1(220) <= to_unsigned(16#86#, 8);
  intdelay_Initial_Val_out_1(221) <= to_unsigned(16#C1#, 8);
  intdelay_Initial_Val_out_1(222) <= to_unsigned(16#1D#, 8);
  intdelay_Initial_Val_out_1(223) <= to_unsigned(16#9E#, 8);
  intdelay_Initial_Val_out_1(224) <= to_unsigned(16#E1#, 8);
  intdelay_Initial_Val_out_1(225) <= to_unsigned(16#F8#, 8);
  intdelay_Initial_Val_out_1(226) <= to_unsigned(16#98#, 8);
  intdelay_Initial_Val_out_1(227) <= to_unsigned(16#11#, 8);
  intdelay_Initial_Val_out_1(228) <= to_unsigned(16#69#, 8);
  intdelay_Initial_Val_out_1(229) <= to_unsigned(16#D9#, 8);
  intdelay_Initial_Val_out_1(230) <= to_unsigned(16#8E#, 8);
  intdelay_Initial_Val_out_1(231) <= to_unsigned(16#94#, 8);
  intdelay_Initial_Val_out_1(232) <= to_unsigned(16#9B#, 8);
  intdelay_Initial_Val_out_1(233) <= to_unsigned(16#1E#, 8);
  intdelay_Initial_Val_out_1(234) <= to_unsigned(16#87#, 8);
  intdelay_Initial_Val_out_1(235) <= to_unsigned(16#E9#, 8);
  intdelay_Initial_Val_out_1(236) <= to_unsigned(16#CE#, 8);
  intdelay_Initial_Val_out_1(237) <= to_unsigned(16#55#, 8);
  intdelay_Initial_Val_out_1(238) <= to_unsigned(16#28#, 8);
  intdelay_Initial_Val_out_1(239) <= to_unsigned(16#DF#, 8);
  intdelay_Initial_Val_out_1(240) <= to_unsigned(16#8C#, 8);
  intdelay_Initial_Val_out_1(241) <= to_unsigned(16#A1#, 8);
  intdelay_Initial_Val_out_1(242) <= to_unsigned(16#89#, 8);
  intdelay_Initial_Val_out_1(243) <= to_unsigned(16#0D#, 8);
  intdelay_Initial_Val_out_1(244) <= to_unsigned(16#BF#, 8);
  intdelay_Initial_Val_out_1(245) <= to_unsigned(16#E6#, 8);
  intdelay_Initial_Val_out_1(246) <= to_unsigned(16#42#, 8);
  intdelay_Initial_Val_out_1(247) <= to_unsigned(16#68#, 8);
  intdelay_Initial_Val_out_1(248) <= to_unsigned(16#41#, 8);
  intdelay_Initial_Val_out_1(249) <= to_unsigned(16#99#, 8);
  intdelay_Initial_Val_out_1(250) <= to_unsigned(16#2D#, 8);
  intdelay_Initial_Val_out_1(251) <= to_unsigned(16#0F#, 8);
  intdelay_Initial_Val_out_1(252) <= to_unsigned(16#B0#, 8);
  intdelay_Initial_Val_out_1(253) <= to_unsigned(16#54#, 8);
  intdelay_Initial_Val_out_1(254) <= to_unsigned(16#BB#, 8);
  intdelay_Initial_Val_out_1(255) <= to_unsigned(16#16#, 8);

  -- #codegen
  intdelay_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_1(0) <= to_unsigned(16#00#, 8);
        intdelay_out_1(1) <= to_unsigned(16#00#, 8);
        intdelay_out_1(2) <= to_unsigned(16#00#, 8);
        intdelay_out_1(3) <= to_unsigned(16#00#, 8);
        intdelay_out_1(4) <= to_unsigned(16#00#, 8);
        intdelay_out_1(5) <= to_unsigned(16#00#, 8);
        intdelay_out_1(6) <= to_unsigned(16#00#, 8);
        intdelay_out_1(7) <= to_unsigned(16#00#, 8);
        intdelay_out_1(8) <= to_unsigned(16#00#, 8);
        intdelay_out_1(9) <= to_unsigned(16#00#, 8);
        intdelay_out_1(10) <= to_unsigned(16#00#, 8);
        intdelay_out_1(11) <= to_unsigned(16#00#, 8);
        intdelay_out_1(12) <= to_unsigned(16#00#, 8);
        intdelay_out_1(13) <= to_unsigned(16#00#, 8);
        intdelay_out_1(14) <= to_unsigned(16#00#, 8);
        intdelay_out_1(15) <= to_unsigned(16#00#, 8);
        intdelay_out_1(16) <= to_unsigned(16#00#, 8);
        intdelay_out_1(17) <= to_unsigned(16#00#, 8);
        intdelay_out_1(18) <= to_unsigned(16#00#, 8);
        intdelay_out_1(19) <= to_unsigned(16#00#, 8);
        intdelay_out_1(20) <= to_unsigned(16#00#, 8);
        intdelay_out_1(21) <= to_unsigned(16#00#, 8);
        intdelay_out_1(22) <= to_unsigned(16#00#, 8);
        intdelay_out_1(23) <= to_unsigned(16#00#, 8);
        intdelay_out_1(24) <= to_unsigned(16#00#, 8);
        intdelay_out_1(25) <= to_unsigned(16#00#, 8);
        intdelay_out_1(26) <= to_unsigned(16#00#, 8);
        intdelay_out_1(27) <= to_unsigned(16#00#, 8);
        intdelay_out_1(28) <= to_unsigned(16#00#, 8);
        intdelay_out_1(29) <= to_unsigned(16#00#, 8);
        intdelay_out_1(30) <= to_unsigned(16#00#, 8);
        intdelay_out_1(31) <= to_unsigned(16#00#, 8);
        intdelay_out_1(32) <= to_unsigned(16#00#, 8);
        intdelay_out_1(33) <= to_unsigned(16#00#, 8);
        intdelay_out_1(34) <= to_unsigned(16#00#, 8);
        intdelay_out_1(35) <= to_unsigned(16#00#, 8);
        intdelay_out_1(36) <= to_unsigned(16#00#, 8);
        intdelay_out_1(37) <= to_unsigned(16#00#, 8);
        intdelay_out_1(38) <= to_unsigned(16#00#, 8);
        intdelay_out_1(39) <= to_unsigned(16#00#, 8);
        intdelay_out_1(40) <= to_unsigned(16#00#, 8);
        intdelay_out_1(41) <= to_unsigned(16#00#, 8);
        intdelay_out_1(42) <= to_unsigned(16#00#, 8);
        intdelay_out_1(43) <= to_unsigned(16#00#, 8);
        intdelay_out_1(44) <= to_unsigned(16#00#, 8);
        intdelay_out_1(45) <= to_unsigned(16#00#, 8);
        intdelay_out_1(46) <= to_unsigned(16#00#, 8);
        intdelay_out_1(47) <= to_unsigned(16#00#, 8);
        intdelay_out_1(48) <= to_unsigned(16#00#, 8);
        intdelay_out_1(49) <= to_unsigned(16#00#, 8);
        intdelay_out_1(50) <= to_unsigned(16#00#, 8);
        intdelay_out_1(51) <= to_unsigned(16#00#, 8);
        intdelay_out_1(52) <= to_unsigned(16#00#, 8);
        intdelay_out_1(53) <= to_unsigned(16#00#, 8);
        intdelay_out_1(54) <= to_unsigned(16#00#, 8);
        intdelay_out_1(55) <= to_unsigned(16#00#, 8);
        intdelay_out_1(56) <= to_unsigned(16#00#, 8);
        intdelay_out_1(57) <= to_unsigned(16#00#, 8);
        intdelay_out_1(58) <= to_unsigned(16#00#, 8);
        intdelay_out_1(59) <= to_unsigned(16#00#, 8);
        intdelay_out_1(60) <= to_unsigned(16#00#, 8);
        intdelay_out_1(61) <= to_unsigned(16#00#, 8);
        intdelay_out_1(62) <= to_unsigned(16#00#, 8);
        intdelay_out_1(63) <= to_unsigned(16#00#, 8);
        intdelay_out_1(64) <= to_unsigned(16#00#, 8);
        intdelay_out_1(65) <= to_unsigned(16#00#, 8);
        intdelay_out_1(66) <= to_unsigned(16#00#, 8);
        intdelay_out_1(67) <= to_unsigned(16#00#, 8);
        intdelay_out_1(68) <= to_unsigned(16#00#, 8);
        intdelay_out_1(69) <= to_unsigned(16#00#, 8);
        intdelay_out_1(70) <= to_unsigned(16#00#, 8);
        intdelay_out_1(71) <= to_unsigned(16#00#, 8);
        intdelay_out_1(72) <= to_unsigned(16#00#, 8);
        intdelay_out_1(73) <= to_unsigned(16#00#, 8);
        intdelay_out_1(74) <= to_unsigned(16#00#, 8);
        intdelay_out_1(75) <= to_unsigned(16#00#, 8);
        intdelay_out_1(76) <= to_unsigned(16#00#, 8);
        intdelay_out_1(77) <= to_unsigned(16#00#, 8);
        intdelay_out_1(78) <= to_unsigned(16#00#, 8);
        intdelay_out_1(79) <= to_unsigned(16#00#, 8);
        intdelay_out_1(80) <= to_unsigned(16#00#, 8);
        intdelay_out_1(81) <= to_unsigned(16#00#, 8);
        intdelay_out_1(82) <= to_unsigned(16#00#, 8);
        intdelay_out_1(83) <= to_unsigned(16#00#, 8);
        intdelay_out_1(84) <= to_unsigned(16#00#, 8);
        intdelay_out_1(85) <= to_unsigned(16#00#, 8);
        intdelay_out_1(86) <= to_unsigned(16#00#, 8);
        intdelay_out_1(87) <= to_unsigned(16#00#, 8);
        intdelay_out_1(88) <= to_unsigned(16#00#, 8);
        intdelay_out_1(89) <= to_unsigned(16#00#, 8);
        intdelay_out_1(90) <= to_unsigned(16#00#, 8);
        intdelay_out_1(91) <= to_unsigned(16#00#, 8);
        intdelay_out_1(92) <= to_unsigned(16#00#, 8);
        intdelay_out_1(93) <= to_unsigned(16#00#, 8);
        intdelay_out_1(94) <= to_unsigned(16#00#, 8);
        intdelay_out_1(95) <= to_unsigned(16#00#, 8);
        intdelay_out_1(96) <= to_unsigned(16#00#, 8);
        intdelay_out_1(97) <= to_unsigned(16#00#, 8);
        intdelay_out_1(98) <= to_unsigned(16#00#, 8);
        intdelay_out_1(99) <= to_unsigned(16#00#, 8);
        intdelay_out_1(100) <= to_unsigned(16#00#, 8);
        intdelay_out_1(101) <= to_unsigned(16#00#, 8);
        intdelay_out_1(102) <= to_unsigned(16#00#, 8);
        intdelay_out_1(103) <= to_unsigned(16#00#, 8);
        intdelay_out_1(104) <= to_unsigned(16#00#, 8);
        intdelay_out_1(105) <= to_unsigned(16#00#, 8);
        intdelay_out_1(106) <= to_unsigned(16#00#, 8);
        intdelay_out_1(107) <= to_unsigned(16#00#, 8);
        intdelay_out_1(108) <= to_unsigned(16#00#, 8);
        intdelay_out_1(109) <= to_unsigned(16#00#, 8);
        intdelay_out_1(110) <= to_unsigned(16#00#, 8);
        intdelay_out_1(111) <= to_unsigned(16#00#, 8);
        intdelay_out_1(112) <= to_unsigned(16#00#, 8);
        intdelay_out_1(113) <= to_unsigned(16#00#, 8);
        intdelay_out_1(114) <= to_unsigned(16#00#, 8);
        intdelay_out_1(115) <= to_unsigned(16#00#, 8);
        intdelay_out_1(116) <= to_unsigned(16#00#, 8);
        intdelay_out_1(117) <= to_unsigned(16#00#, 8);
        intdelay_out_1(118) <= to_unsigned(16#00#, 8);
        intdelay_out_1(119) <= to_unsigned(16#00#, 8);
        intdelay_out_1(120) <= to_unsigned(16#00#, 8);
        intdelay_out_1(121) <= to_unsigned(16#00#, 8);
        intdelay_out_1(122) <= to_unsigned(16#00#, 8);
        intdelay_out_1(123) <= to_unsigned(16#00#, 8);
        intdelay_out_1(124) <= to_unsigned(16#00#, 8);
        intdelay_out_1(125) <= to_unsigned(16#00#, 8);
        intdelay_out_1(126) <= to_unsigned(16#00#, 8);
        intdelay_out_1(127) <= to_unsigned(16#00#, 8);
        intdelay_out_1(128) <= to_unsigned(16#00#, 8);
        intdelay_out_1(129) <= to_unsigned(16#00#, 8);
        intdelay_out_1(130) <= to_unsigned(16#00#, 8);
        intdelay_out_1(131) <= to_unsigned(16#00#, 8);
        intdelay_out_1(132) <= to_unsigned(16#00#, 8);
        intdelay_out_1(133) <= to_unsigned(16#00#, 8);
        intdelay_out_1(134) <= to_unsigned(16#00#, 8);
        intdelay_out_1(135) <= to_unsigned(16#00#, 8);
        intdelay_out_1(136) <= to_unsigned(16#00#, 8);
        intdelay_out_1(137) <= to_unsigned(16#00#, 8);
        intdelay_out_1(138) <= to_unsigned(16#00#, 8);
        intdelay_out_1(139) <= to_unsigned(16#00#, 8);
        intdelay_out_1(140) <= to_unsigned(16#00#, 8);
        intdelay_out_1(141) <= to_unsigned(16#00#, 8);
        intdelay_out_1(142) <= to_unsigned(16#00#, 8);
        intdelay_out_1(143) <= to_unsigned(16#00#, 8);
        intdelay_out_1(144) <= to_unsigned(16#00#, 8);
        intdelay_out_1(145) <= to_unsigned(16#00#, 8);
        intdelay_out_1(146) <= to_unsigned(16#00#, 8);
        intdelay_out_1(147) <= to_unsigned(16#00#, 8);
        intdelay_out_1(148) <= to_unsigned(16#00#, 8);
        intdelay_out_1(149) <= to_unsigned(16#00#, 8);
        intdelay_out_1(150) <= to_unsigned(16#00#, 8);
        intdelay_out_1(151) <= to_unsigned(16#00#, 8);
        intdelay_out_1(152) <= to_unsigned(16#00#, 8);
        intdelay_out_1(153) <= to_unsigned(16#00#, 8);
        intdelay_out_1(154) <= to_unsigned(16#00#, 8);
        intdelay_out_1(155) <= to_unsigned(16#00#, 8);
        intdelay_out_1(156) <= to_unsigned(16#00#, 8);
        intdelay_out_1(157) <= to_unsigned(16#00#, 8);
        intdelay_out_1(158) <= to_unsigned(16#00#, 8);
        intdelay_out_1(159) <= to_unsigned(16#00#, 8);
        intdelay_out_1(160) <= to_unsigned(16#00#, 8);
        intdelay_out_1(161) <= to_unsigned(16#00#, 8);
        intdelay_out_1(162) <= to_unsigned(16#00#, 8);
        intdelay_out_1(163) <= to_unsigned(16#00#, 8);
        intdelay_out_1(164) <= to_unsigned(16#00#, 8);
        intdelay_out_1(165) <= to_unsigned(16#00#, 8);
        intdelay_out_1(166) <= to_unsigned(16#00#, 8);
        intdelay_out_1(167) <= to_unsigned(16#00#, 8);
        intdelay_out_1(168) <= to_unsigned(16#00#, 8);
        intdelay_out_1(169) <= to_unsigned(16#00#, 8);
        intdelay_out_1(170) <= to_unsigned(16#00#, 8);
        intdelay_out_1(171) <= to_unsigned(16#00#, 8);
        intdelay_out_1(172) <= to_unsigned(16#00#, 8);
        intdelay_out_1(173) <= to_unsigned(16#00#, 8);
        intdelay_out_1(174) <= to_unsigned(16#00#, 8);
        intdelay_out_1(175) <= to_unsigned(16#00#, 8);
        intdelay_out_1(176) <= to_unsigned(16#00#, 8);
        intdelay_out_1(177) <= to_unsigned(16#00#, 8);
        intdelay_out_1(178) <= to_unsigned(16#00#, 8);
        intdelay_out_1(179) <= to_unsigned(16#00#, 8);
        intdelay_out_1(180) <= to_unsigned(16#00#, 8);
        intdelay_out_1(181) <= to_unsigned(16#00#, 8);
        intdelay_out_1(182) <= to_unsigned(16#00#, 8);
        intdelay_out_1(183) <= to_unsigned(16#00#, 8);
        intdelay_out_1(184) <= to_unsigned(16#00#, 8);
        intdelay_out_1(185) <= to_unsigned(16#00#, 8);
        intdelay_out_1(186) <= to_unsigned(16#00#, 8);
        intdelay_out_1(187) <= to_unsigned(16#00#, 8);
        intdelay_out_1(188) <= to_unsigned(16#00#, 8);
        intdelay_out_1(189) <= to_unsigned(16#00#, 8);
        intdelay_out_1(190) <= to_unsigned(16#00#, 8);
        intdelay_out_1(191) <= to_unsigned(16#00#, 8);
        intdelay_out_1(192) <= to_unsigned(16#00#, 8);
        intdelay_out_1(193) <= to_unsigned(16#00#, 8);
        intdelay_out_1(194) <= to_unsigned(16#00#, 8);
        intdelay_out_1(195) <= to_unsigned(16#00#, 8);
        intdelay_out_1(196) <= to_unsigned(16#00#, 8);
        intdelay_out_1(197) <= to_unsigned(16#00#, 8);
        intdelay_out_1(198) <= to_unsigned(16#00#, 8);
        intdelay_out_1(199) <= to_unsigned(16#00#, 8);
        intdelay_out_1(200) <= to_unsigned(16#00#, 8);
        intdelay_out_1(201) <= to_unsigned(16#00#, 8);
        intdelay_out_1(202) <= to_unsigned(16#00#, 8);
        intdelay_out_1(203) <= to_unsigned(16#00#, 8);
        intdelay_out_1(204) <= to_unsigned(16#00#, 8);
        intdelay_out_1(205) <= to_unsigned(16#00#, 8);
        intdelay_out_1(206) <= to_unsigned(16#00#, 8);
        intdelay_out_1(207) <= to_unsigned(16#00#, 8);
        intdelay_out_1(208) <= to_unsigned(16#00#, 8);
        intdelay_out_1(209) <= to_unsigned(16#00#, 8);
        intdelay_out_1(210) <= to_unsigned(16#00#, 8);
        intdelay_out_1(211) <= to_unsigned(16#00#, 8);
        intdelay_out_1(212) <= to_unsigned(16#00#, 8);
        intdelay_out_1(213) <= to_unsigned(16#00#, 8);
        intdelay_out_1(214) <= to_unsigned(16#00#, 8);
        intdelay_out_1(215) <= to_unsigned(16#00#, 8);
        intdelay_out_1(216) <= to_unsigned(16#00#, 8);
        intdelay_out_1(217) <= to_unsigned(16#00#, 8);
        intdelay_out_1(218) <= to_unsigned(16#00#, 8);
        intdelay_out_1(219) <= to_unsigned(16#00#, 8);
        intdelay_out_1(220) <= to_unsigned(16#00#, 8);
        intdelay_out_1(221) <= to_unsigned(16#00#, 8);
        intdelay_out_1(222) <= to_unsigned(16#00#, 8);
        intdelay_out_1(223) <= to_unsigned(16#00#, 8);
        intdelay_out_1(224) <= to_unsigned(16#00#, 8);
        intdelay_out_1(225) <= to_unsigned(16#00#, 8);
        intdelay_out_1(226) <= to_unsigned(16#00#, 8);
        intdelay_out_1(227) <= to_unsigned(16#00#, 8);
        intdelay_out_1(228) <= to_unsigned(16#00#, 8);
        intdelay_out_1(229) <= to_unsigned(16#00#, 8);
        intdelay_out_1(230) <= to_unsigned(16#00#, 8);
        intdelay_out_1(231) <= to_unsigned(16#00#, 8);
        intdelay_out_1(232) <= to_unsigned(16#00#, 8);
        intdelay_out_1(233) <= to_unsigned(16#00#, 8);
        intdelay_out_1(234) <= to_unsigned(16#00#, 8);
        intdelay_out_1(235) <= to_unsigned(16#00#, 8);
        intdelay_out_1(236) <= to_unsigned(16#00#, 8);
        intdelay_out_1(237) <= to_unsigned(16#00#, 8);
        intdelay_out_1(238) <= to_unsigned(16#00#, 8);
        intdelay_out_1(239) <= to_unsigned(16#00#, 8);
        intdelay_out_1(240) <= to_unsigned(16#00#, 8);
        intdelay_out_1(241) <= to_unsigned(16#00#, 8);
        intdelay_out_1(242) <= to_unsigned(16#00#, 8);
        intdelay_out_1(243) <= to_unsigned(16#00#, 8);
        intdelay_out_1(244) <= to_unsigned(16#00#, 8);
        intdelay_out_1(245) <= to_unsigned(16#00#, 8);
        intdelay_out_1(246) <= to_unsigned(16#00#, 8);
        intdelay_out_1(247) <= to_unsigned(16#00#, 8);
        intdelay_out_1(248) <= to_unsigned(16#00#, 8);
        intdelay_out_1(249) <= to_unsigned(16#00#, 8);
        intdelay_out_1(250) <= to_unsigned(16#00#, 8);
        intdelay_out_1(251) <= to_unsigned(16#00#, 8);
        intdelay_out_1(252) <= to_unsigned(16#00#, 8);
        intdelay_out_1(253) <= to_unsigned(16#00#, 8);
        intdelay_out_1(254) <= to_unsigned(16#00#, 8);
        intdelay_out_1(255) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_1(0) <= sbox(0);
        intdelay_out_1(1) <= sbox(1);
        intdelay_out_1(2) <= sbox(2);
        intdelay_out_1(3) <= sbox(3);
        intdelay_out_1(4) <= sbox(4);
        intdelay_out_1(5) <= sbox(5);
        intdelay_out_1(6) <= sbox(6);
        intdelay_out_1(7) <= sbox(7);
        intdelay_out_1(8) <= sbox(8);
        intdelay_out_1(9) <= sbox(9);
        intdelay_out_1(10) <= sbox(10);
        intdelay_out_1(11) <= sbox(11);
        intdelay_out_1(12) <= sbox(12);
        intdelay_out_1(13) <= sbox(13);
        intdelay_out_1(14) <= sbox(14);
        intdelay_out_1(15) <= sbox(15);
        intdelay_out_1(16) <= sbox(16);
        intdelay_out_1(17) <= sbox(17);
        intdelay_out_1(18) <= sbox(18);
        intdelay_out_1(19) <= sbox(19);
        intdelay_out_1(20) <= sbox(20);
        intdelay_out_1(21) <= sbox(21);
        intdelay_out_1(22) <= sbox(22);
        intdelay_out_1(23) <= sbox(23);
        intdelay_out_1(24) <= sbox(24);
        intdelay_out_1(25) <= sbox(25);
        intdelay_out_1(26) <= sbox(26);
        intdelay_out_1(27) <= sbox(27);
        intdelay_out_1(28) <= sbox(28);
        intdelay_out_1(29) <= sbox(29);
        intdelay_out_1(30) <= sbox(30);
        intdelay_out_1(31) <= sbox(31);
        intdelay_out_1(32) <= sbox(32);
        intdelay_out_1(33) <= sbox(33);
        intdelay_out_1(34) <= sbox(34);
        intdelay_out_1(35) <= sbox(35);
        intdelay_out_1(36) <= sbox(36);
        intdelay_out_1(37) <= sbox(37);
        intdelay_out_1(38) <= sbox(38);
        intdelay_out_1(39) <= sbox(39);
        intdelay_out_1(40) <= sbox(40);
        intdelay_out_1(41) <= sbox(41);
        intdelay_out_1(42) <= sbox(42);
        intdelay_out_1(43) <= sbox(43);
        intdelay_out_1(44) <= sbox(44);
        intdelay_out_1(45) <= sbox(45);
        intdelay_out_1(46) <= sbox(46);
        intdelay_out_1(47) <= sbox(47);
        intdelay_out_1(48) <= sbox(48);
        intdelay_out_1(49) <= sbox(49);
        intdelay_out_1(50) <= sbox(50);
        intdelay_out_1(51) <= sbox(51);
        intdelay_out_1(52) <= sbox(52);
        intdelay_out_1(53) <= sbox(53);
        intdelay_out_1(54) <= sbox(54);
        intdelay_out_1(55) <= sbox(55);
        intdelay_out_1(56) <= sbox(56);
        intdelay_out_1(57) <= sbox(57);
        intdelay_out_1(58) <= sbox(58);
        intdelay_out_1(59) <= sbox(59);
        intdelay_out_1(60) <= sbox(60);
        intdelay_out_1(61) <= sbox(61);
        intdelay_out_1(62) <= sbox(62);
        intdelay_out_1(63) <= sbox(63);
        intdelay_out_1(64) <= sbox(64);
        intdelay_out_1(65) <= sbox(65);
        intdelay_out_1(66) <= sbox(66);
        intdelay_out_1(67) <= sbox(67);
        intdelay_out_1(68) <= sbox(68);
        intdelay_out_1(69) <= sbox(69);
        intdelay_out_1(70) <= sbox(70);
        intdelay_out_1(71) <= sbox(71);
        intdelay_out_1(72) <= sbox(72);
        intdelay_out_1(73) <= sbox(73);
        intdelay_out_1(74) <= sbox(74);
        intdelay_out_1(75) <= sbox(75);
        intdelay_out_1(76) <= sbox(76);
        intdelay_out_1(77) <= sbox(77);
        intdelay_out_1(78) <= sbox(78);
        intdelay_out_1(79) <= sbox(79);
        intdelay_out_1(80) <= sbox(80);
        intdelay_out_1(81) <= sbox(81);
        intdelay_out_1(82) <= sbox(82);
        intdelay_out_1(83) <= sbox(83);
        intdelay_out_1(84) <= sbox(84);
        intdelay_out_1(85) <= sbox(85);
        intdelay_out_1(86) <= sbox(86);
        intdelay_out_1(87) <= sbox(87);
        intdelay_out_1(88) <= sbox(88);
        intdelay_out_1(89) <= sbox(89);
        intdelay_out_1(90) <= sbox(90);
        intdelay_out_1(91) <= sbox(91);
        intdelay_out_1(92) <= sbox(92);
        intdelay_out_1(93) <= sbox(93);
        intdelay_out_1(94) <= sbox(94);
        intdelay_out_1(95) <= sbox(95);
        intdelay_out_1(96) <= sbox(96);
        intdelay_out_1(97) <= sbox(97);
        intdelay_out_1(98) <= sbox(98);
        intdelay_out_1(99) <= sbox(99);
        intdelay_out_1(100) <= sbox(100);
        intdelay_out_1(101) <= sbox(101);
        intdelay_out_1(102) <= sbox(102);
        intdelay_out_1(103) <= sbox(103);
        intdelay_out_1(104) <= sbox(104);
        intdelay_out_1(105) <= sbox(105);
        intdelay_out_1(106) <= sbox(106);
        intdelay_out_1(107) <= sbox(107);
        intdelay_out_1(108) <= sbox(108);
        intdelay_out_1(109) <= sbox(109);
        intdelay_out_1(110) <= sbox(110);
        intdelay_out_1(111) <= sbox(111);
        intdelay_out_1(112) <= sbox(112);
        intdelay_out_1(113) <= sbox(113);
        intdelay_out_1(114) <= sbox(114);
        intdelay_out_1(115) <= sbox(115);
        intdelay_out_1(116) <= sbox(116);
        intdelay_out_1(117) <= sbox(117);
        intdelay_out_1(118) <= sbox(118);
        intdelay_out_1(119) <= sbox(119);
        intdelay_out_1(120) <= sbox(120);
        intdelay_out_1(121) <= sbox(121);
        intdelay_out_1(122) <= sbox(122);
        intdelay_out_1(123) <= sbox(123);
        intdelay_out_1(124) <= sbox(124);
        intdelay_out_1(125) <= sbox(125);
        intdelay_out_1(126) <= sbox(126);
        intdelay_out_1(127) <= sbox(127);
        intdelay_out_1(128) <= sbox(128);
        intdelay_out_1(129) <= sbox(129);
        intdelay_out_1(130) <= sbox(130);
        intdelay_out_1(131) <= sbox(131);
        intdelay_out_1(132) <= sbox(132);
        intdelay_out_1(133) <= sbox(133);
        intdelay_out_1(134) <= sbox(134);
        intdelay_out_1(135) <= sbox(135);
        intdelay_out_1(136) <= sbox(136);
        intdelay_out_1(137) <= sbox(137);
        intdelay_out_1(138) <= sbox(138);
        intdelay_out_1(139) <= sbox(139);
        intdelay_out_1(140) <= sbox(140);
        intdelay_out_1(141) <= sbox(141);
        intdelay_out_1(142) <= sbox(142);
        intdelay_out_1(143) <= sbox(143);
        intdelay_out_1(144) <= sbox(144);
        intdelay_out_1(145) <= sbox(145);
        intdelay_out_1(146) <= sbox(146);
        intdelay_out_1(147) <= sbox(147);
        intdelay_out_1(148) <= sbox(148);
        intdelay_out_1(149) <= sbox(149);
        intdelay_out_1(150) <= sbox(150);
        intdelay_out_1(151) <= sbox(151);
        intdelay_out_1(152) <= sbox(152);
        intdelay_out_1(153) <= sbox(153);
        intdelay_out_1(154) <= sbox(154);
        intdelay_out_1(155) <= sbox(155);
        intdelay_out_1(156) <= sbox(156);
        intdelay_out_1(157) <= sbox(157);
        intdelay_out_1(158) <= sbox(158);
        intdelay_out_1(159) <= sbox(159);
        intdelay_out_1(160) <= sbox(160);
        intdelay_out_1(161) <= sbox(161);
        intdelay_out_1(162) <= sbox(162);
        intdelay_out_1(163) <= sbox(163);
        intdelay_out_1(164) <= sbox(164);
        intdelay_out_1(165) <= sbox(165);
        intdelay_out_1(166) <= sbox(166);
        intdelay_out_1(167) <= sbox(167);
        intdelay_out_1(168) <= sbox(168);
        intdelay_out_1(169) <= sbox(169);
        intdelay_out_1(170) <= sbox(170);
        intdelay_out_1(171) <= sbox(171);
        intdelay_out_1(172) <= sbox(172);
        intdelay_out_1(173) <= sbox(173);
        intdelay_out_1(174) <= sbox(174);
        intdelay_out_1(175) <= sbox(175);
        intdelay_out_1(176) <= sbox(176);
        intdelay_out_1(177) <= sbox(177);
        intdelay_out_1(178) <= sbox(178);
        intdelay_out_1(179) <= sbox(179);
        intdelay_out_1(180) <= sbox(180);
        intdelay_out_1(181) <= sbox(181);
        intdelay_out_1(182) <= sbox(182);
        intdelay_out_1(183) <= sbox(183);
        intdelay_out_1(184) <= sbox(184);
        intdelay_out_1(185) <= sbox(185);
        intdelay_out_1(186) <= sbox(186);
        intdelay_out_1(187) <= sbox(187);
        intdelay_out_1(188) <= sbox(188);
        intdelay_out_1(189) <= sbox(189);
        intdelay_out_1(190) <= sbox(190);
        intdelay_out_1(191) <= sbox(191);
        intdelay_out_1(192) <= sbox(192);
        intdelay_out_1(193) <= sbox(193);
        intdelay_out_1(194) <= sbox(194);
        intdelay_out_1(195) <= sbox(195);
        intdelay_out_1(196) <= sbox(196);
        intdelay_out_1(197) <= sbox(197);
        intdelay_out_1(198) <= sbox(198);
        intdelay_out_1(199) <= sbox(199);
        intdelay_out_1(200) <= sbox(200);
        intdelay_out_1(201) <= sbox(201);
        intdelay_out_1(202) <= sbox(202);
        intdelay_out_1(203) <= sbox(203);
        intdelay_out_1(204) <= sbox(204);
        intdelay_out_1(205) <= sbox(205);
        intdelay_out_1(206) <= sbox(206);
        intdelay_out_1(207) <= sbox(207);
        intdelay_out_1(208) <= sbox(208);
        intdelay_out_1(209) <= sbox(209);
        intdelay_out_1(210) <= sbox(210);
        intdelay_out_1(211) <= sbox(211);
        intdelay_out_1(212) <= sbox(212);
        intdelay_out_1(213) <= sbox(213);
        intdelay_out_1(214) <= sbox(214);
        intdelay_out_1(215) <= sbox(215);
        intdelay_out_1(216) <= sbox(216);
        intdelay_out_1(217) <= sbox(217);
        intdelay_out_1(218) <= sbox(218);
        intdelay_out_1(219) <= sbox(219);
        intdelay_out_1(220) <= sbox(220);
        intdelay_out_1(221) <= sbox(221);
        intdelay_out_1(222) <= sbox(222);
        intdelay_out_1(223) <= sbox(223);
        intdelay_out_1(224) <= sbox(224);
        intdelay_out_1(225) <= sbox(225);
        intdelay_out_1(226) <= sbox(226);
        intdelay_out_1(227) <= sbox(227);
        intdelay_out_1(228) <= sbox(228);
        intdelay_out_1(229) <= sbox(229);
        intdelay_out_1(230) <= sbox(230);
        intdelay_out_1(231) <= sbox(231);
        intdelay_out_1(232) <= sbox(232);
        intdelay_out_1(233) <= sbox(233);
        intdelay_out_1(234) <= sbox(234);
        intdelay_out_1(235) <= sbox(235);
        intdelay_out_1(236) <= sbox(236);
        intdelay_out_1(237) <= sbox(237);
        intdelay_out_1(238) <= sbox(238);
        intdelay_out_1(239) <= sbox(239);
        intdelay_out_1(240) <= sbox(240);
        intdelay_out_1(241) <= sbox(241);
        intdelay_out_1(242) <= sbox(242);
        intdelay_out_1(243) <= sbox(243);
        intdelay_out_1(244) <= sbox(244);
        intdelay_out_1(245) <= sbox(245);
        intdelay_out_1(246) <= sbox(246);
        intdelay_out_1(247) <= sbox(247);
        intdelay_out_1(248) <= sbox(248);
        intdelay_out_1(249) <= sbox(249);
        intdelay_out_1(250) <= sbox(250);
        intdelay_out_1(251) <= sbox(251);
        intdelay_out_1(252) <= sbox(252);
        intdelay_out_1(253) <= sbox(253);
        intdelay_out_1(254) <= sbox(254);
        intdelay_out_1(255) <= sbox(255);
      END IF;
    END IF;
  END PROCESS intdelay_process;


  
  sbox(0) <= intdelay_Initial_Val_out_1(0) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(0);
  
  sbox(1) <= intdelay_Initial_Val_out_1(1) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(1);
  
  sbox(2) <= intdelay_Initial_Val_out_1(2) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(2);
  
  sbox(3) <= intdelay_Initial_Val_out_1(3) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(3);
  
  sbox(4) <= intdelay_Initial_Val_out_1(4) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(4);
  
  sbox(5) <= intdelay_Initial_Val_out_1(5) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(5);
  
  sbox(6) <= intdelay_Initial_Val_out_1(6) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(6);
  
  sbox(7) <= intdelay_Initial_Val_out_1(7) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(7);
  
  sbox(8) <= intdelay_Initial_Val_out_1(8) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(8);
  
  sbox(9) <= intdelay_Initial_Val_out_1(9) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(9);
  
  sbox(10) <= intdelay_Initial_Val_out_1(10) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(10);
  
  sbox(11) <= intdelay_Initial_Val_out_1(11) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(11);
  
  sbox(12) <= intdelay_Initial_Val_out_1(12) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(12);
  
  sbox(13) <= intdelay_Initial_Val_out_1(13) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(13);
  
  sbox(14) <= intdelay_Initial_Val_out_1(14) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(14);
  
  sbox(15) <= intdelay_Initial_Val_out_1(15) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(15);
  
  sbox(16) <= intdelay_Initial_Val_out_1(16) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(16);
  
  sbox(17) <= intdelay_Initial_Val_out_1(17) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(17);
  
  sbox(18) <= intdelay_Initial_Val_out_1(18) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(18);
  
  sbox(19) <= intdelay_Initial_Val_out_1(19) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(19);
  
  sbox(20) <= intdelay_Initial_Val_out_1(20) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(20);
  
  sbox(21) <= intdelay_Initial_Val_out_1(21) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(21);
  
  sbox(22) <= intdelay_Initial_Val_out_1(22) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(22);
  
  sbox(23) <= intdelay_Initial_Val_out_1(23) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(23);
  
  sbox(24) <= intdelay_Initial_Val_out_1(24) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(24);
  
  sbox(25) <= intdelay_Initial_Val_out_1(25) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(25);
  
  sbox(26) <= intdelay_Initial_Val_out_1(26) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(26);
  
  sbox(27) <= intdelay_Initial_Val_out_1(27) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(27);
  
  sbox(28) <= intdelay_Initial_Val_out_1(28) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(28);
  
  sbox(29) <= intdelay_Initial_Val_out_1(29) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(29);
  
  sbox(30) <= intdelay_Initial_Val_out_1(30) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(30);
  
  sbox(31) <= intdelay_Initial_Val_out_1(31) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(31);
  
  sbox(32) <= intdelay_Initial_Val_out_1(32) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(32);
  
  sbox(33) <= intdelay_Initial_Val_out_1(33) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(33);
  
  sbox(34) <= intdelay_Initial_Val_out_1(34) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(34);
  
  sbox(35) <= intdelay_Initial_Val_out_1(35) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(35);
  
  sbox(36) <= intdelay_Initial_Val_out_1(36) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(36);
  
  sbox(37) <= intdelay_Initial_Val_out_1(37) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(37);
  
  sbox(38) <= intdelay_Initial_Val_out_1(38) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(38);
  
  sbox(39) <= intdelay_Initial_Val_out_1(39) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(39);
  
  sbox(40) <= intdelay_Initial_Val_out_1(40) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(40);
  
  sbox(41) <= intdelay_Initial_Val_out_1(41) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(41);
  
  sbox(42) <= intdelay_Initial_Val_out_1(42) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(42);
  
  sbox(43) <= intdelay_Initial_Val_out_1(43) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(43);
  
  sbox(44) <= intdelay_Initial_Val_out_1(44) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(44);
  
  sbox(45) <= intdelay_Initial_Val_out_1(45) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(45);
  
  sbox(46) <= intdelay_Initial_Val_out_1(46) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(46);
  
  sbox(47) <= intdelay_Initial_Val_out_1(47) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(47);
  
  sbox(48) <= intdelay_Initial_Val_out_1(48) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(48);
  
  sbox(49) <= intdelay_Initial_Val_out_1(49) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(49);
  
  sbox(50) <= intdelay_Initial_Val_out_1(50) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(50);
  
  sbox(51) <= intdelay_Initial_Val_out_1(51) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(51);
  
  sbox(52) <= intdelay_Initial_Val_out_1(52) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(52);
  
  sbox(53) <= intdelay_Initial_Val_out_1(53) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(53);
  
  sbox(54) <= intdelay_Initial_Val_out_1(54) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(54);
  
  sbox(55) <= intdelay_Initial_Val_out_1(55) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(55);
  
  sbox(56) <= intdelay_Initial_Val_out_1(56) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(56);
  
  sbox(57) <= intdelay_Initial_Val_out_1(57) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(57);
  
  sbox(58) <= intdelay_Initial_Val_out_1(58) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(58);
  
  sbox(59) <= intdelay_Initial_Val_out_1(59) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(59);
  
  sbox(60) <= intdelay_Initial_Val_out_1(60) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(60);
  
  sbox(61) <= intdelay_Initial_Val_out_1(61) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(61);
  
  sbox(62) <= intdelay_Initial_Val_out_1(62) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(62);
  
  sbox(63) <= intdelay_Initial_Val_out_1(63) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(63);
  
  sbox(64) <= intdelay_Initial_Val_out_1(64) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(64);
  
  sbox(65) <= intdelay_Initial_Val_out_1(65) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(65);
  
  sbox(66) <= intdelay_Initial_Val_out_1(66) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(66);
  
  sbox(67) <= intdelay_Initial_Val_out_1(67) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(67);
  
  sbox(68) <= intdelay_Initial_Val_out_1(68) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(68);
  
  sbox(69) <= intdelay_Initial_Val_out_1(69) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(69);
  
  sbox(70) <= intdelay_Initial_Val_out_1(70) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(70);
  
  sbox(71) <= intdelay_Initial_Val_out_1(71) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(71);
  
  sbox(72) <= intdelay_Initial_Val_out_1(72) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(72);
  
  sbox(73) <= intdelay_Initial_Val_out_1(73) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(73);
  
  sbox(74) <= intdelay_Initial_Val_out_1(74) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(74);
  
  sbox(75) <= intdelay_Initial_Val_out_1(75) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(75);
  
  sbox(76) <= intdelay_Initial_Val_out_1(76) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(76);
  
  sbox(77) <= intdelay_Initial_Val_out_1(77) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(77);
  
  sbox(78) <= intdelay_Initial_Val_out_1(78) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(78);
  
  sbox(79) <= intdelay_Initial_Val_out_1(79) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(79);
  
  sbox(80) <= intdelay_Initial_Val_out_1(80) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(80);
  
  sbox(81) <= intdelay_Initial_Val_out_1(81) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(81);
  
  sbox(82) <= intdelay_Initial_Val_out_1(82) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(82);
  
  sbox(83) <= intdelay_Initial_Val_out_1(83) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(83);
  
  sbox(84) <= intdelay_Initial_Val_out_1(84) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(84);
  
  sbox(85) <= intdelay_Initial_Val_out_1(85) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(85);
  
  sbox(86) <= intdelay_Initial_Val_out_1(86) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(86);
  
  sbox(87) <= intdelay_Initial_Val_out_1(87) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(87);
  
  sbox(88) <= intdelay_Initial_Val_out_1(88) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(88);
  
  sbox(89) <= intdelay_Initial_Val_out_1(89) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(89);
  
  sbox(90) <= intdelay_Initial_Val_out_1(90) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(90);
  
  sbox(91) <= intdelay_Initial_Val_out_1(91) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(91);
  
  sbox(92) <= intdelay_Initial_Val_out_1(92) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(92);
  
  sbox(93) <= intdelay_Initial_Val_out_1(93) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(93);
  
  sbox(94) <= intdelay_Initial_Val_out_1(94) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(94);
  
  sbox(95) <= intdelay_Initial_Val_out_1(95) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(95);
  
  sbox(96) <= intdelay_Initial_Val_out_1(96) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(96);
  
  sbox(97) <= intdelay_Initial_Val_out_1(97) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(97);
  
  sbox(98) <= intdelay_Initial_Val_out_1(98) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(98);
  
  sbox(99) <= intdelay_Initial_Val_out_1(99) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(99);
  
  sbox(100) <= intdelay_Initial_Val_out_1(100) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(100);
  
  sbox(101) <= intdelay_Initial_Val_out_1(101) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(101);
  
  sbox(102) <= intdelay_Initial_Val_out_1(102) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(102);
  
  sbox(103) <= intdelay_Initial_Val_out_1(103) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(103);
  
  sbox(104) <= intdelay_Initial_Val_out_1(104) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(104);
  
  sbox(105) <= intdelay_Initial_Val_out_1(105) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(105);
  
  sbox(106) <= intdelay_Initial_Val_out_1(106) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(106);
  
  sbox(107) <= intdelay_Initial_Val_out_1(107) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(107);
  
  sbox(108) <= intdelay_Initial_Val_out_1(108) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(108);
  
  sbox(109) <= intdelay_Initial_Val_out_1(109) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(109);
  
  sbox(110) <= intdelay_Initial_Val_out_1(110) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(110);
  
  sbox(111) <= intdelay_Initial_Val_out_1(111) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(111);
  
  sbox(112) <= intdelay_Initial_Val_out_1(112) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(112);
  
  sbox(113) <= intdelay_Initial_Val_out_1(113) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(113);
  
  sbox(114) <= intdelay_Initial_Val_out_1(114) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(114);
  
  sbox(115) <= intdelay_Initial_Val_out_1(115) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(115);
  
  sbox(116) <= intdelay_Initial_Val_out_1(116) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(116);
  
  sbox(117) <= intdelay_Initial_Val_out_1(117) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(117);
  
  sbox(118) <= intdelay_Initial_Val_out_1(118) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(118);
  
  sbox(119) <= intdelay_Initial_Val_out_1(119) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(119);
  
  sbox(120) <= intdelay_Initial_Val_out_1(120) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(120);
  
  sbox(121) <= intdelay_Initial_Val_out_1(121) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(121);
  
  sbox(122) <= intdelay_Initial_Val_out_1(122) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(122);
  
  sbox(123) <= intdelay_Initial_Val_out_1(123) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(123);
  
  sbox(124) <= intdelay_Initial_Val_out_1(124) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(124);
  
  sbox(125) <= intdelay_Initial_Val_out_1(125) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(125);
  
  sbox(126) <= intdelay_Initial_Val_out_1(126) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(126);
  
  sbox(127) <= intdelay_Initial_Val_out_1(127) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(127);
  
  sbox(128) <= intdelay_Initial_Val_out_1(128) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(128);
  
  sbox(129) <= intdelay_Initial_Val_out_1(129) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(129);
  
  sbox(130) <= intdelay_Initial_Val_out_1(130) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(130);
  
  sbox(131) <= intdelay_Initial_Val_out_1(131) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(131);
  
  sbox(132) <= intdelay_Initial_Val_out_1(132) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(132);
  
  sbox(133) <= intdelay_Initial_Val_out_1(133) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(133);
  
  sbox(134) <= intdelay_Initial_Val_out_1(134) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(134);
  
  sbox(135) <= intdelay_Initial_Val_out_1(135) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(135);
  
  sbox(136) <= intdelay_Initial_Val_out_1(136) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(136);
  
  sbox(137) <= intdelay_Initial_Val_out_1(137) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(137);
  
  sbox(138) <= intdelay_Initial_Val_out_1(138) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(138);
  
  sbox(139) <= intdelay_Initial_Val_out_1(139) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(139);
  
  sbox(140) <= intdelay_Initial_Val_out_1(140) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(140);
  
  sbox(141) <= intdelay_Initial_Val_out_1(141) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(141);
  
  sbox(142) <= intdelay_Initial_Val_out_1(142) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(142);
  
  sbox(143) <= intdelay_Initial_Val_out_1(143) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(143);
  
  sbox(144) <= intdelay_Initial_Val_out_1(144) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(144);
  
  sbox(145) <= intdelay_Initial_Val_out_1(145) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(145);
  
  sbox(146) <= intdelay_Initial_Val_out_1(146) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(146);
  
  sbox(147) <= intdelay_Initial_Val_out_1(147) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(147);
  
  sbox(148) <= intdelay_Initial_Val_out_1(148) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(148);
  
  sbox(149) <= intdelay_Initial_Val_out_1(149) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(149);
  
  sbox(150) <= intdelay_Initial_Val_out_1(150) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(150);
  
  sbox(151) <= intdelay_Initial_Val_out_1(151) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(151);
  
  sbox(152) <= intdelay_Initial_Val_out_1(152) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(152);
  
  sbox(153) <= intdelay_Initial_Val_out_1(153) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(153);
  
  sbox(154) <= intdelay_Initial_Val_out_1(154) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(154);
  
  sbox(155) <= intdelay_Initial_Val_out_1(155) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(155);
  
  sbox(156) <= intdelay_Initial_Val_out_1(156) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(156);
  
  sbox(157) <= intdelay_Initial_Val_out_1(157) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(157);
  
  sbox(158) <= intdelay_Initial_Val_out_1(158) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(158);
  
  sbox(159) <= intdelay_Initial_Val_out_1(159) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(159);
  
  sbox(160) <= intdelay_Initial_Val_out_1(160) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(160);
  
  sbox(161) <= intdelay_Initial_Val_out_1(161) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(161);
  
  sbox(162) <= intdelay_Initial_Val_out_1(162) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(162);
  
  sbox(163) <= intdelay_Initial_Val_out_1(163) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(163);
  
  sbox(164) <= intdelay_Initial_Val_out_1(164) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(164);
  
  sbox(165) <= intdelay_Initial_Val_out_1(165) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(165);
  
  sbox(166) <= intdelay_Initial_Val_out_1(166) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(166);
  
  sbox(167) <= intdelay_Initial_Val_out_1(167) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(167);
  
  sbox(168) <= intdelay_Initial_Val_out_1(168) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(168);
  
  sbox(169) <= intdelay_Initial_Val_out_1(169) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(169);
  
  sbox(170) <= intdelay_Initial_Val_out_1(170) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(170);
  
  sbox(171) <= intdelay_Initial_Val_out_1(171) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(171);
  
  sbox(172) <= intdelay_Initial_Val_out_1(172) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(172);
  
  sbox(173) <= intdelay_Initial_Val_out_1(173) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(173);
  
  sbox(174) <= intdelay_Initial_Val_out_1(174) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(174);
  
  sbox(175) <= intdelay_Initial_Val_out_1(175) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(175);
  
  sbox(176) <= intdelay_Initial_Val_out_1(176) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(176);
  
  sbox(177) <= intdelay_Initial_Val_out_1(177) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(177);
  
  sbox(178) <= intdelay_Initial_Val_out_1(178) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(178);
  
  sbox(179) <= intdelay_Initial_Val_out_1(179) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(179);
  
  sbox(180) <= intdelay_Initial_Val_out_1(180) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(180);
  
  sbox(181) <= intdelay_Initial_Val_out_1(181) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(181);
  
  sbox(182) <= intdelay_Initial_Val_out_1(182) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(182);
  
  sbox(183) <= intdelay_Initial_Val_out_1(183) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(183);
  
  sbox(184) <= intdelay_Initial_Val_out_1(184) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(184);
  
  sbox(185) <= intdelay_Initial_Val_out_1(185) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(185);
  
  sbox(186) <= intdelay_Initial_Val_out_1(186) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(186);
  
  sbox(187) <= intdelay_Initial_Val_out_1(187) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(187);
  
  sbox(188) <= intdelay_Initial_Val_out_1(188) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(188);
  
  sbox(189) <= intdelay_Initial_Val_out_1(189) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(189);
  
  sbox(190) <= intdelay_Initial_Val_out_1(190) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(190);
  
  sbox(191) <= intdelay_Initial_Val_out_1(191) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(191);
  
  sbox(192) <= intdelay_Initial_Val_out_1(192) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(192);
  
  sbox(193) <= intdelay_Initial_Val_out_1(193) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(193);
  
  sbox(194) <= intdelay_Initial_Val_out_1(194) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(194);
  
  sbox(195) <= intdelay_Initial_Val_out_1(195) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(195);
  
  sbox(196) <= intdelay_Initial_Val_out_1(196) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(196);
  
  sbox(197) <= intdelay_Initial_Val_out_1(197) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(197);
  
  sbox(198) <= intdelay_Initial_Val_out_1(198) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(198);
  
  sbox(199) <= intdelay_Initial_Val_out_1(199) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(199);
  
  sbox(200) <= intdelay_Initial_Val_out_1(200) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(200);
  
  sbox(201) <= intdelay_Initial_Val_out_1(201) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(201);
  
  sbox(202) <= intdelay_Initial_Val_out_1(202) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(202);
  
  sbox(203) <= intdelay_Initial_Val_out_1(203) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(203);
  
  sbox(204) <= intdelay_Initial_Val_out_1(204) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(204);
  
  sbox(205) <= intdelay_Initial_Val_out_1(205) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(205);
  
  sbox(206) <= intdelay_Initial_Val_out_1(206) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(206);
  
  sbox(207) <= intdelay_Initial_Val_out_1(207) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(207);
  
  sbox(208) <= intdelay_Initial_Val_out_1(208) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(208);
  
  sbox(209) <= intdelay_Initial_Val_out_1(209) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(209);
  
  sbox(210) <= intdelay_Initial_Val_out_1(210) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(210);
  
  sbox(211) <= intdelay_Initial_Val_out_1(211) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(211);
  
  sbox(212) <= intdelay_Initial_Val_out_1(212) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(212);
  
  sbox(213) <= intdelay_Initial_Val_out_1(213) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(213);
  
  sbox(214) <= intdelay_Initial_Val_out_1(214) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(214);
  
  sbox(215) <= intdelay_Initial_Val_out_1(215) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(215);
  
  sbox(216) <= intdelay_Initial_Val_out_1(216) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(216);
  
  sbox(217) <= intdelay_Initial_Val_out_1(217) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(217);
  
  sbox(218) <= intdelay_Initial_Val_out_1(218) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(218);
  
  sbox(219) <= intdelay_Initial_Val_out_1(219) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(219);
  
  sbox(220) <= intdelay_Initial_Val_out_1(220) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(220);
  
  sbox(221) <= intdelay_Initial_Val_out_1(221) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(221);
  
  sbox(222) <= intdelay_Initial_Val_out_1(222) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(222);
  
  sbox(223) <= intdelay_Initial_Val_out_1(223) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(223);
  
  sbox(224) <= intdelay_Initial_Val_out_1(224) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(224);
  
  sbox(225) <= intdelay_Initial_Val_out_1(225) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(225);
  
  sbox(226) <= intdelay_Initial_Val_out_1(226) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(226);
  
  sbox(227) <= intdelay_Initial_Val_out_1(227) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(227);
  
  sbox(228) <= intdelay_Initial_Val_out_1(228) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(228);
  
  sbox(229) <= intdelay_Initial_Val_out_1(229) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(229);
  
  sbox(230) <= intdelay_Initial_Val_out_1(230) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(230);
  
  sbox(231) <= intdelay_Initial_Val_out_1(231) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(231);
  
  sbox(232) <= intdelay_Initial_Val_out_1(232) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(232);
  
  sbox(233) <= intdelay_Initial_Val_out_1(233) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(233);
  
  sbox(234) <= intdelay_Initial_Val_out_1(234) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(234);
  
  sbox(235) <= intdelay_Initial_Val_out_1(235) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(235);
  
  sbox(236) <= intdelay_Initial_Val_out_1(236) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(236);
  
  sbox(237) <= intdelay_Initial_Val_out_1(237) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(237);
  
  sbox(238) <= intdelay_Initial_Val_out_1(238) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(238);
  
  sbox(239) <= intdelay_Initial_Val_out_1(239) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(239);
  
  sbox(240) <= intdelay_Initial_Val_out_1(240) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(240);
  
  sbox(241) <= intdelay_Initial_Val_out_1(241) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(241);
  
  sbox(242) <= intdelay_Initial_Val_out_1(242) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(242);
  
  sbox(243) <= intdelay_Initial_Val_out_1(243) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(243);
  
  sbox(244) <= intdelay_Initial_Val_out_1(244) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(244);
  
  sbox(245) <= intdelay_Initial_Val_out_1(245) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(245);
  
  sbox(246) <= intdelay_Initial_Val_out_1(246) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(246);
  
  sbox(247) <= intdelay_Initial_Val_out_1(247) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(247);
  
  sbox(248) <= intdelay_Initial_Val_out_1(248) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(248);
  
  sbox(249) <= intdelay_Initial_Val_out_1(249) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(249);
  
  sbox(250) <= intdelay_Initial_Val_out_1(250) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(250);
  
  sbox(251) <= intdelay_Initial_Val_out_1(251) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(251);
  
  sbox(252) <= intdelay_Initial_Val_out_1(252) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(252);
  
  sbox(253) <= intdelay_Initial_Val_out_1(253) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(253);
  
  sbox(254) <= intdelay_Initial_Val_out_1(254) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(254);
  
  sbox(255) <= intdelay_Initial_Val_out_1(255) WHEN intdelay_ctrl_delay_out_1 = '0' ELSE
      intdelay_out_1(255);

  const_expression_14 <= to_unsigned(16#0001#, 16);

  jj <= ii_4 sll 2;

  const_expression_15 <= to_unsigned(16#04#, 8);

  out0_55 <= jj - const_expression_15;

  iii <= to_unsigned(16#01#, 8);

  out0_56 <= out0_55 + iii;

  intdelay_ctrl_const_out_2 <= '1';

  intdelay_ctrl_delay1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_ctrl_delay_out_2 <= '0';
      ELSIF enb = '1' THEN
        intdelay_ctrl_delay_out_2 <= intdelay_ctrl_const_out_2;
      END IF;
    END IF;
  END PROCESS intdelay_ctrl_delay1_process;


  intdelay_Initial_Val_out_2(0) <= to_unsigned(16#01#, 8);
  intdelay_Initial_Val_out_2(1) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(2) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(3) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(4) <= to_unsigned(16#02#, 8);
  intdelay_Initial_Val_out_2(5) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(6) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(7) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(8) <= to_unsigned(16#04#, 8);
  intdelay_Initial_Val_out_2(9) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(10) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(11) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(12) <= to_unsigned(16#08#, 8);
  intdelay_Initial_Val_out_2(13) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(14) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(15) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(16) <= to_unsigned(16#10#, 8);
  intdelay_Initial_Val_out_2(17) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(18) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(19) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(20) <= to_unsigned(16#20#, 8);
  intdelay_Initial_Val_out_2(21) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(22) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(23) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(24) <= to_unsigned(16#40#, 8);
  intdelay_Initial_Val_out_2(25) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(26) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(27) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(28) <= to_unsigned(16#80#, 8);
  intdelay_Initial_Val_out_2(29) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(30) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(31) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(32) <= to_unsigned(16#1B#, 8);
  intdelay_Initial_Val_out_2(33) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(34) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(35) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(36) <= to_unsigned(16#36#, 8);
  intdelay_Initial_Val_out_2(37) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(38) <= to_unsigned(16#00#, 8);
  intdelay_Initial_Val_out_2(39) <= to_unsigned(16#00#, 8);

  intdelay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        intdelay_out_2(0) <= to_unsigned(16#00#, 8);
        intdelay_out_2(1) <= to_unsigned(16#00#, 8);
        intdelay_out_2(2) <= to_unsigned(16#00#, 8);
        intdelay_out_2(3) <= to_unsigned(16#00#, 8);
        intdelay_out_2(4) <= to_unsigned(16#00#, 8);
        intdelay_out_2(5) <= to_unsigned(16#00#, 8);
        intdelay_out_2(6) <= to_unsigned(16#00#, 8);
        intdelay_out_2(7) <= to_unsigned(16#00#, 8);
        intdelay_out_2(8) <= to_unsigned(16#00#, 8);
        intdelay_out_2(9) <= to_unsigned(16#00#, 8);
        intdelay_out_2(10) <= to_unsigned(16#00#, 8);
        intdelay_out_2(11) <= to_unsigned(16#00#, 8);
        intdelay_out_2(12) <= to_unsigned(16#00#, 8);
        intdelay_out_2(13) <= to_unsigned(16#00#, 8);
        intdelay_out_2(14) <= to_unsigned(16#00#, 8);
        intdelay_out_2(15) <= to_unsigned(16#00#, 8);
        intdelay_out_2(16) <= to_unsigned(16#00#, 8);
        intdelay_out_2(17) <= to_unsigned(16#00#, 8);
        intdelay_out_2(18) <= to_unsigned(16#00#, 8);
        intdelay_out_2(19) <= to_unsigned(16#00#, 8);
        intdelay_out_2(20) <= to_unsigned(16#00#, 8);
        intdelay_out_2(21) <= to_unsigned(16#00#, 8);
        intdelay_out_2(22) <= to_unsigned(16#00#, 8);
        intdelay_out_2(23) <= to_unsigned(16#00#, 8);
        intdelay_out_2(24) <= to_unsigned(16#00#, 8);
        intdelay_out_2(25) <= to_unsigned(16#00#, 8);
        intdelay_out_2(26) <= to_unsigned(16#00#, 8);
        intdelay_out_2(27) <= to_unsigned(16#00#, 8);
        intdelay_out_2(28) <= to_unsigned(16#00#, 8);
        intdelay_out_2(29) <= to_unsigned(16#00#, 8);
        intdelay_out_2(30) <= to_unsigned(16#00#, 8);
        intdelay_out_2(31) <= to_unsigned(16#00#, 8);
        intdelay_out_2(32) <= to_unsigned(16#00#, 8);
        intdelay_out_2(33) <= to_unsigned(16#00#, 8);
        intdelay_out_2(34) <= to_unsigned(16#00#, 8);
        intdelay_out_2(35) <= to_unsigned(16#00#, 8);
        intdelay_out_2(36) <= to_unsigned(16#00#, 8);
        intdelay_out_2(37) <= to_unsigned(16#00#, 8);
        intdelay_out_2(38) <= to_unsigned(16#00#, 8);
        intdelay_out_2(39) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        intdelay_out_2(0) <= Rcon(0);
        intdelay_out_2(1) <= Rcon(1);
        intdelay_out_2(2) <= Rcon(2);
        intdelay_out_2(3) <= Rcon(3);
        intdelay_out_2(4) <= Rcon(4);
        intdelay_out_2(5) <= Rcon(5);
        intdelay_out_2(6) <= Rcon(6);
        intdelay_out_2(7) <= Rcon(7);
        intdelay_out_2(8) <= Rcon(8);
        intdelay_out_2(9) <= Rcon(9);
        intdelay_out_2(10) <= Rcon(10);
        intdelay_out_2(11) <= Rcon(11);
        intdelay_out_2(12) <= Rcon(12);
        intdelay_out_2(13) <= Rcon(13);
        intdelay_out_2(14) <= Rcon(14);
        intdelay_out_2(15) <= Rcon(15);
        intdelay_out_2(16) <= Rcon(16);
        intdelay_out_2(17) <= Rcon(17);
        intdelay_out_2(18) <= Rcon(18);
        intdelay_out_2(19) <= Rcon(19);
        intdelay_out_2(20) <= Rcon(20);
        intdelay_out_2(21) <= Rcon(21);
        intdelay_out_2(22) <= Rcon(22);
        intdelay_out_2(23) <= Rcon(23);
        intdelay_out_2(24) <= Rcon(24);
        intdelay_out_2(25) <= Rcon(25);
        intdelay_out_2(26) <= Rcon(26);
        intdelay_out_2(27) <= Rcon(27);
        intdelay_out_2(28) <= Rcon(28);
        intdelay_out_2(29) <= Rcon(29);
        intdelay_out_2(30) <= Rcon(30);
        intdelay_out_2(31) <= Rcon(31);
        intdelay_out_2(32) <= Rcon(32);
        intdelay_out_2(33) <= Rcon(33);
        intdelay_out_2(34) <= Rcon(34);
        intdelay_out_2(35) <= Rcon(35);
        intdelay_out_2(36) <= Rcon(36);
        intdelay_out_2(37) <= Rcon(37);
        intdelay_out_2(38) <= Rcon(38);
        intdelay_out_2(39) <= Rcon(39);
      END IF;
    END IF;
  END PROCESS intdelay2_process;


  
  Rcon(0) <= intdelay_Initial_Val_out_2(0) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(0);
  
  Rcon(1) <= intdelay_Initial_Val_out_2(1) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(1);
  
  Rcon(2) <= intdelay_Initial_Val_out_2(2) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(2);
  
  Rcon(3) <= intdelay_Initial_Val_out_2(3) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(3);
  
  Rcon(4) <= intdelay_Initial_Val_out_2(4) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(4);
  
  Rcon(5) <= intdelay_Initial_Val_out_2(5) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(5);
  
  Rcon(6) <= intdelay_Initial_Val_out_2(6) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(6);
  
  Rcon(7) <= intdelay_Initial_Val_out_2(7) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(7);
  
  Rcon(8) <= intdelay_Initial_Val_out_2(8) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(8);
  
  Rcon(9) <= intdelay_Initial_Val_out_2(9) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(9);
  
  Rcon(10) <= intdelay_Initial_Val_out_2(10) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(10);
  
  Rcon(11) <= intdelay_Initial_Val_out_2(11) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(11);
  
  Rcon(12) <= intdelay_Initial_Val_out_2(12) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(12);
  
  Rcon(13) <= intdelay_Initial_Val_out_2(13) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(13);
  
  Rcon(14) <= intdelay_Initial_Val_out_2(14) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(14);
  
  Rcon(15) <= intdelay_Initial_Val_out_2(15) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(15);
  
  Rcon(16) <= intdelay_Initial_Val_out_2(16) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(16);
  
  Rcon(17) <= intdelay_Initial_Val_out_2(17) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(17);
  
  Rcon(18) <= intdelay_Initial_Val_out_2(18) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(18);
  
  Rcon(19) <= intdelay_Initial_Val_out_2(19) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(19);
  
  Rcon(20) <= intdelay_Initial_Val_out_2(20) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(20);
  
  Rcon(21) <= intdelay_Initial_Val_out_2(21) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(21);
  
  Rcon(22) <= intdelay_Initial_Val_out_2(22) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(22);
  
  Rcon(23) <= intdelay_Initial_Val_out_2(23) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(23);
  
  Rcon(24) <= intdelay_Initial_Val_out_2(24) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(24);
  
  Rcon(25) <= intdelay_Initial_Val_out_2(25) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(25);
  
  Rcon(26) <= intdelay_Initial_Val_out_2(26) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(26);
  
  Rcon(27) <= intdelay_Initial_Val_out_2(27) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(27);
  
  Rcon(28) <= intdelay_Initial_Val_out_2(28) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(28);
  
  Rcon(29) <= intdelay_Initial_Val_out_2(29) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(29);
  
  Rcon(30) <= intdelay_Initial_Val_out_2(30) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(30);
  
  Rcon(31) <= intdelay_Initial_Val_out_2(31) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(31);
  
  Rcon(32) <= intdelay_Initial_Val_out_2(32) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(32);
  
  Rcon(33) <= intdelay_Initial_Val_out_2(33) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(33);
  
  Rcon(34) <= intdelay_Initial_Val_out_2(34) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(34);
  
  Rcon(35) <= intdelay_Initial_Val_out_2(35) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(35);
  
  Rcon(36) <= intdelay_Initial_Val_out_2(36) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(36);
  
  Rcon(37) <= intdelay_Initial_Val_out_2(37) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(37);
  
  Rcon(38) <= intdelay_Initial_Val_out_2(38) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(38);
  
  Rcon(39) <= intdelay_Initial_Val_out_2(39) WHEN intdelay_ctrl_delay_out_2 = '0' ELSE
      intdelay_out_2(39);

  
  out0_57 <= Rcon(0) WHEN out0_56 = to_unsigned(16#01#, 8) ELSE
      Rcon(1) WHEN out0_56 = to_unsigned(16#02#, 8) ELSE
      Rcon(2) WHEN out0_56 = to_unsigned(16#03#, 8) ELSE
      Rcon(3) WHEN out0_56 = to_unsigned(16#04#, 8) ELSE
      Rcon(4) WHEN out0_56 = to_unsigned(16#05#, 8) ELSE
      Rcon(5) WHEN out0_56 = to_unsigned(16#06#, 8) ELSE
      Rcon(6) WHEN out0_56 = to_unsigned(16#07#, 8) ELSE
      Rcon(7) WHEN out0_56 = to_unsigned(16#08#, 8) ELSE
      Rcon(8) WHEN out0_56 = to_unsigned(16#09#, 8) ELSE
      Rcon(9) WHEN out0_56 = to_unsigned(16#0A#, 8) ELSE
      Rcon(10) WHEN out0_56 = to_unsigned(16#0B#, 8) ELSE
      Rcon(11) WHEN out0_56 = to_unsigned(16#0C#, 8) ELSE
      Rcon(12) WHEN out0_56 = to_unsigned(16#0D#, 8) ELSE
      Rcon(13) WHEN out0_56 = to_unsigned(16#0E#, 8) ELSE
      Rcon(14) WHEN out0_56 = to_unsigned(16#0F#, 8) ELSE
      Rcon(15) WHEN out0_56 = to_unsigned(16#10#, 8) ELSE
      Rcon(16) WHEN out0_56 = to_unsigned(16#11#, 8) ELSE
      Rcon(17) WHEN out0_56 = to_unsigned(16#12#, 8) ELSE
      Rcon(18) WHEN out0_56 = to_unsigned(16#13#, 8) ELSE
      Rcon(19) WHEN out0_56 = to_unsigned(16#14#, 8) ELSE
      Rcon(20) WHEN out0_56 = to_unsigned(16#15#, 8) ELSE
      Rcon(21) WHEN out0_56 = to_unsigned(16#16#, 8) ELSE
      Rcon(22) WHEN out0_56 = to_unsigned(16#17#, 8) ELSE
      Rcon(23) WHEN out0_56 = to_unsigned(16#18#, 8) ELSE
      Rcon(24) WHEN out0_56 = to_unsigned(16#19#, 8) ELSE
      Rcon(25) WHEN out0_56 = to_unsigned(16#1A#, 8) ELSE
      Rcon(26) WHEN out0_56 = to_unsigned(16#1B#, 8) ELSE
      Rcon(27) WHEN out0_56 = to_unsigned(16#1C#, 8) ELSE
      Rcon(28) WHEN out0_56 = to_unsigned(16#1D#, 8) ELSE
      Rcon(29) WHEN out0_56 = to_unsigned(16#1E#, 8) ELSE
      Rcon(30) WHEN out0_56 = to_unsigned(16#1F#, 8) ELSE
      Rcon(31) WHEN out0_56 = to_unsigned(16#20#, 8) ELSE
      Rcon(32) WHEN out0_56 = to_unsigned(16#21#, 8) ELSE
      Rcon(33) WHEN out0_56 = to_unsigned(16#22#, 8) ELSE
      Rcon(34) WHEN out0_56 = to_unsigned(16#23#, 8) ELSE
      Rcon(35) WHEN out0_56 = to_unsigned(16#24#, 8) ELSE
      Rcon(36) WHEN out0_56 = to_unsigned(16#25#, 8) ELSE
      Rcon(37) WHEN out0_56 = to_unsigned(16#26#, 8) ELSE
      Rcon(38) WHEN out0_56 = to_unsigned(16#27#, 8) ELSE
      Rcon(39);

  const_expression_16 <= to_unsigned(16#04#, 8);

  out0_58 <= jj - const_expression_16;

  iii_1 <= to_unsigned(16#02#, 8);

  out0_59 <= out0_58 + iii_1;

  
  out0_60 <= Rcon(0) WHEN out0_59 = to_unsigned(16#01#, 8) ELSE
      Rcon(1) WHEN out0_59 = to_unsigned(16#02#, 8) ELSE
      Rcon(2) WHEN out0_59 = to_unsigned(16#03#, 8) ELSE
      Rcon(3) WHEN out0_59 = to_unsigned(16#04#, 8) ELSE
      Rcon(4) WHEN out0_59 = to_unsigned(16#05#, 8) ELSE
      Rcon(5) WHEN out0_59 = to_unsigned(16#06#, 8) ELSE
      Rcon(6) WHEN out0_59 = to_unsigned(16#07#, 8) ELSE
      Rcon(7) WHEN out0_59 = to_unsigned(16#08#, 8) ELSE
      Rcon(8) WHEN out0_59 = to_unsigned(16#09#, 8) ELSE
      Rcon(9) WHEN out0_59 = to_unsigned(16#0A#, 8) ELSE
      Rcon(10) WHEN out0_59 = to_unsigned(16#0B#, 8) ELSE
      Rcon(11) WHEN out0_59 = to_unsigned(16#0C#, 8) ELSE
      Rcon(12) WHEN out0_59 = to_unsigned(16#0D#, 8) ELSE
      Rcon(13) WHEN out0_59 = to_unsigned(16#0E#, 8) ELSE
      Rcon(14) WHEN out0_59 = to_unsigned(16#0F#, 8) ELSE
      Rcon(15) WHEN out0_59 = to_unsigned(16#10#, 8) ELSE
      Rcon(16) WHEN out0_59 = to_unsigned(16#11#, 8) ELSE
      Rcon(17) WHEN out0_59 = to_unsigned(16#12#, 8) ELSE
      Rcon(18) WHEN out0_59 = to_unsigned(16#13#, 8) ELSE
      Rcon(19) WHEN out0_59 = to_unsigned(16#14#, 8) ELSE
      Rcon(20) WHEN out0_59 = to_unsigned(16#15#, 8) ELSE
      Rcon(21) WHEN out0_59 = to_unsigned(16#16#, 8) ELSE
      Rcon(22) WHEN out0_59 = to_unsigned(16#17#, 8) ELSE
      Rcon(23) WHEN out0_59 = to_unsigned(16#18#, 8) ELSE
      Rcon(24) WHEN out0_59 = to_unsigned(16#19#, 8) ELSE
      Rcon(25) WHEN out0_59 = to_unsigned(16#1A#, 8) ELSE
      Rcon(26) WHEN out0_59 = to_unsigned(16#1B#, 8) ELSE
      Rcon(27) WHEN out0_59 = to_unsigned(16#1C#, 8) ELSE
      Rcon(28) WHEN out0_59 = to_unsigned(16#1D#, 8) ELSE
      Rcon(29) WHEN out0_59 = to_unsigned(16#1E#, 8) ELSE
      Rcon(30) WHEN out0_59 = to_unsigned(16#1F#, 8) ELSE
      Rcon(31) WHEN out0_59 = to_unsigned(16#20#, 8) ELSE
      Rcon(32) WHEN out0_59 = to_unsigned(16#21#, 8) ELSE
      Rcon(33) WHEN out0_59 = to_unsigned(16#22#, 8) ELSE
      Rcon(34) WHEN out0_59 = to_unsigned(16#23#, 8) ELSE
      Rcon(35) WHEN out0_59 = to_unsigned(16#24#, 8) ELSE
      Rcon(36) WHEN out0_59 = to_unsigned(16#25#, 8) ELSE
      Rcon(37) WHEN out0_59 = to_unsigned(16#26#, 8) ELSE
      Rcon(38) WHEN out0_59 = to_unsigned(16#27#, 8) ELSE
      Rcon(39);

  const_expression_17 <= to_unsigned(16#04#, 8);

  out0_61 <= jj - const_expression_17;

  iii_2 <= to_unsigned(16#03#, 8);

  out0_62 <= out0_61 + iii_2;

  
  out0_63 <= Rcon(0) WHEN out0_62 = to_unsigned(16#01#, 8) ELSE
      Rcon(1) WHEN out0_62 = to_unsigned(16#02#, 8) ELSE
      Rcon(2) WHEN out0_62 = to_unsigned(16#03#, 8) ELSE
      Rcon(3) WHEN out0_62 = to_unsigned(16#04#, 8) ELSE
      Rcon(4) WHEN out0_62 = to_unsigned(16#05#, 8) ELSE
      Rcon(5) WHEN out0_62 = to_unsigned(16#06#, 8) ELSE
      Rcon(6) WHEN out0_62 = to_unsigned(16#07#, 8) ELSE
      Rcon(7) WHEN out0_62 = to_unsigned(16#08#, 8) ELSE
      Rcon(8) WHEN out0_62 = to_unsigned(16#09#, 8) ELSE
      Rcon(9) WHEN out0_62 = to_unsigned(16#0A#, 8) ELSE
      Rcon(10) WHEN out0_62 = to_unsigned(16#0B#, 8) ELSE
      Rcon(11) WHEN out0_62 = to_unsigned(16#0C#, 8) ELSE
      Rcon(12) WHEN out0_62 = to_unsigned(16#0D#, 8) ELSE
      Rcon(13) WHEN out0_62 = to_unsigned(16#0E#, 8) ELSE
      Rcon(14) WHEN out0_62 = to_unsigned(16#0F#, 8) ELSE
      Rcon(15) WHEN out0_62 = to_unsigned(16#10#, 8) ELSE
      Rcon(16) WHEN out0_62 = to_unsigned(16#11#, 8) ELSE
      Rcon(17) WHEN out0_62 = to_unsigned(16#12#, 8) ELSE
      Rcon(18) WHEN out0_62 = to_unsigned(16#13#, 8) ELSE
      Rcon(19) WHEN out0_62 = to_unsigned(16#14#, 8) ELSE
      Rcon(20) WHEN out0_62 = to_unsigned(16#15#, 8) ELSE
      Rcon(21) WHEN out0_62 = to_unsigned(16#16#, 8) ELSE
      Rcon(22) WHEN out0_62 = to_unsigned(16#17#, 8) ELSE
      Rcon(23) WHEN out0_62 = to_unsigned(16#18#, 8) ELSE
      Rcon(24) WHEN out0_62 = to_unsigned(16#19#, 8) ELSE
      Rcon(25) WHEN out0_62 = to_unsigned(16#1A#, 8) ELSE
      Rcon(26) WHEN out0_62 = to_unsigned(16#1B#, 8) ELSE
      Rcon(27) WHEN out0_62 = to_unsigned(16#1C#, 8) ELSE
      Rcon(28) WHEN out0_62 = to_unsigned(16#1D#, 8) ELSE
      Rcon(29) WHEN out0_62 = to_unsigned(16#1E#, 8) ELSE
      Rcon(30) WHEN out0_62 = to_unsigned(16#1F#, 8) ELSE
      Rcon(31) WHEN out0_62 = to_unsigned(16#20#, 8) ELSE
      Rcon(32) WHEN out0_62 = to_unsigned(16#21#, 8) ELSE
      Rcon(33) WHEN out0_62 = to_unsigned(16#22#, 8) ELSE
      Rcon(34) WHEN out0_62 = to_unsigned(16#23#, 8) ELSE
      Rcon(35) WHEN out0_62 = to_unsigned(16#24#, 8) ELSE
      Rcon(36) WHEN out0_62 = to_unsigned(16#25#, 8) ELSE
      Rcon(37) WHEN out0_62 = to_unsigned(16#26#, 8) ELSE
      Rcon(38) WHEN out0_62 = to_unsigned(16#27#, 8) ELSE
      Rcon(39);

  const_expression_18 <= to_unsigned(16#04#, 8);

  out0_64 <= jj - const_expression_18;

  iii_3 <= to_unsigned(16#04#, 8);

  out0_65 <= out0_64 + iii_3;

  
  out0_66 <= Rcon(0) WHEN out0_65 = to_unsigned(16#01#, 8) ELSE
      Rcon(1) WHEN out0_65 = to_unsigned(16#02#, 8) ELSE
      Rcon(2) WHEN out0_65 = to_unsigned(16#03#, 8) ELSE
      Rcon(3) WHEN out0_65 = to_unsigned(16#04#, 8) ELSE
      Rcon(4) WHEN out0_65 = to_unsigned(16#05#, 8) ELSE
      Rcon(5) WHEN out0_65 = to_unsigned(16#06#, 8) ELSE
      Rcon(6) WHEN out0_65 = to_unsigned(16#07#, 8) ELSE
      Rcon(7) WHEN out0_65 = to_unsigned(16#08#, 8) ELSE
      Rcon(8) WHEN out0_65 = to_unsigned(16#09#, 8) ELSE
      Rcon(9) WHEN out0_65 = to_unsigned(16#0A#, 8) ELSE
      Rcon(10) WHEN out0_65 = to_unsigned(16#0B#, 8) ELSE
      Rcon(11) WHEN out0_65 = to_unsigned(16#0C#, 8) ELSE
      Rcon(12) WHEN out0_65 = to_unsigned(16#0D#, 8) ELSE
      Rcon(13) WHEN out0_65 = to_unsigned(16#0E#, 8) ELSE
      Rcon(14) WHEN out0_65 = to_unsigned(16#0F#, 8) ELSE
      Rcon(15) WHEN out0_65 = to_unsigned(16#10#, 8) ELSE
      Rcon(16) WHEN out0_65 = to_unsigned(16#11#, 8) ELSE
      Rcon(17) WHEN out0_65 = to_unsigned(16#12#, 8) ELSE
      Rcon(18) WHEN out0_65 = to_unsigned(16#13#, 8) ELSE
      Rcon(19) WHEN out0_65 = to_unsigned(16#14#, 8) ELSE
      Rcon(20) WHEN out0_65 = to_unsigned(16#15#, 8) ELSE
      Rcon(21) WHEN out0_65 = to_unsigned(16#16#, 8) ELSE
      Rcon(22) WHEN out0_65 = to_unsigned(16#17#, 8) ELSE
      Rcon(23) WHEN out0_65 = to_unsigned(16#18#, 8) ELSE
      Rcon(24) WHEN out0_65 = to_unsigned(16#19#, 8) ELSE
      Rcon(25) WHEN out0_65 = to_unsigned(16#1A#, 8) ELSE
      Rcon(26) WHEN out0_65 = to_unsigned(16#1B#, 8) ELSE
      Rcon(27) WHEN out0_65 = to_unsigned(16#1C#, 8) ELSE
      Rcon(28) WHEN out0_65 = to_unsigned(16#1D#, 8) ELSE
      Rcon(29) WHEN out0_65 = to_unsigned(16#1E#, 8) ELSE
      Rcon(30) WHEN out0_65 = to_unsigned(16#1F#, 8) ELSE
      Rcon(31) WHEN out0_65 = to_unsigned(16#20#, 8) ELSE
      Rcon(32) WHEN out0_65 = to_unsigned(16#21#, 8) ELSE
      Rcon(33) WHEN out0_65 = to_unsigned(16#22#, 8) ELSE
      Rcon(34) WHEN out0_65 = to_unsigned(16#23#, 8) ELSE
      Rcon(35) WHEN out0_65 = to_unsigned(16#24#, 8) ELSE
      Rcon(36) WHEN out0_65 = to_unsigned(16#25#, 8) ELSE
      Rcon(37) WHEN out0_65 = to_unsigned(16#26#, 8) ELSE
      Rcon(38) WHEN out0_65 = to_unsigned(16#27#, 8) ELSE
      Rcon(39);

  
  out0_67(0) <= k2(0) WHEN out0_5 = '0' ELSE
      k2(0);
  
  out0_67(1) <= k2(1) WHEN out0_5 = '0' ELSE
      k2(1);
  
  out0_67(2) <= k2(2) WHEN out0_5 = '0' ELSE
      k2(2);
  
  out0_67(3) <= k2(3) WHEN out0_5 = '0' ELSE
      k2(3);

  
  k2_2(0) <= out0_67(0) WHEN out0_9 = '0' ELSE
      k2_1(0);
  
  k2_2(1) <= out0_67(1) WHEN out0_9 = '0' ELSE
      k2_1(1);
  
  k2_2(2) <= out0_67(2) WHEN out0_9 = '0' ELSE
      k2_1(2);
  
  k2_2(3) <= out0_67(3) WHEN out0_9 = '0' ELSE
      k2_1(3);

  
  out0_68(0) <= k2(0) WHEN out0_10 = '0' ELSE
      k2(0);
  
  out0_68(1) <= k2(1) WHEN out0_10 = '0' ELSE
      k2(1);
  
  out0_68(2) <= k2(2) WHEN out0_10 = '0' ELSE
      k2(2);
  
  out0_68(3) <= k2(3) WHEN out0_10 = '0' ELSE
      k2(3);

  
  out0_69(0) <= out0_68(0) WHEN out0_12 = '0' ELSE
      k2(0);
  
  out0_69(1) <= out0_68(1) WHEN out0_12 = '0' ELSE
      k2(1);
  
  out0_69(2) <= out0_68(2) WHEN out0_12 = '0' ELSE
      k2(2);
  
  out0_69(3) <= out0_68(3) WHEN out0_12 = '0' ELSE
      k2(3);

  
  out0_70(0) <= out0_69(0) WHEN out0_14 = '0' ELSE
      k2(0);
  
  out0_70(1) <= out0_69(1) WHEN out0_14 = '0' ELSE
      k2(1);
  
  out0_70(2) <= out0_69(2) WHEN out0_14 = '0' ELSE
      k2(2);
  
  out0_70(3) <= out0_69(3) WHEN out0_14 = '0' ELSE
      k2(3);

  
  out0_71(0) <= out0_70(0) WHEN out0_16 = '0' ELSE
      k2(0);
  
  out0_71(1) <= out0_70(1) WHEN out0_16 = '0' ELSE
      k2(1);
  
  out0_71(2) <= out0_70(2) WHEN out0_16 = '0' ELSE
      k2(2);
  
  out0_71(3) <= out0_70(3) WHEN out0_16 = '0' ELSE
      k2(3);

  
  out0_72(0) <= out0_71(0) WHEN out0_18 = '0' ELSE
      k2(0);
  
  out0_72(1) <= out0_71(1) WHEN out0_18 = '0' ELSE
      k2(1);
  
  out0_72(2) <= out0_71(2) WHEN out0_18 = '0' ELSE
      k2(2);
  
  out0_72(3) <= out0_71(3) WHEN out0_18 = '0' ELSE
      k2(3);

  
  out0_73(0) <= out0_72(0) WHEN out0_20 = '0' ELSE
      k2(0);
  
  out0_73(1) <= out0_72(1) WHEN out0_20 = '0' ELSE
      k2(1);
  
  out0_73(2) <= out0_72(2) WHEN out0_20 = '0' ELSE
      k2(2);
  
  out0_73(3) <= out0_72(3) WHEN out0_20 = '0' ELSE
      k2(3);

  
  out0_74(0) <= out0_73(0) WHEN out0_22 = '0' ELSE
      k2_2(0);
  
  out0_74(1) <= out0_73(1) WHEN out0_22 = '0' ELSE
      k2_2(1);
  
  out0_74(2) <= out0_73(2) WHEN out0_22 = '0' ELSE
      k2_2(2);
  
  out0_74(3) <= out0_73(3) WHEN out0_22 = '0' ELSE
      k2_2(3);

  
  k2_3(0) <= out0_74(0) WHEN out0_24 = '0' ELSE
      k2(0);
  
  k2_3(1) <= out0_74(1) WHEN out0_24 = '0' ELSE
      k2(1);
  
  k2_3(2) <= out0_74(2) WHEN out0_24 = '0' ELSE
      k2(2);
  
  k2_3(3) <= out0_74(3) WHEN out0_24 = '0' ELSE
      k2(3);

  intdelay10_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        k2(0) <= to_unsigned(16#00#, 8);
        k2(1) <= to_unsigned(16#00#, 8);
        k2(2) <= to_unsigned(16#00#, 8);
        k2(3) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        k2(0) <= k2_3(0);
        k2(1) <= k2_3(1);
        k2(2) <= k2_3(2);
        k2(3) <= k2_3(3);
      END IF;
    END IF;
  END PROCESS intdelay10_process;


  k2_4(0) <= out0_57;
  k2_4(1) <= k2(1);
  k2_4(2) <= k2(2);
  k2_4(3) <= k2(3);

  k2_5(0) <= k2_4(0);
  k2_5(1) <= out0_60;
  k2_5(2) <= k2_4(2);
  k2_5(3) <= k2_4(3);

  k2_6(0) <= k2_5(0);
  k2_6(1) <= k2_5(1);
  k2_6(2) <= out0_63;
  k2_6(3) <= k2_5(3);

  k2_1(0) <= k2_6(0);
  k2_1(1) <= k2_6(1);
  k2_1(2) <= k2_6(2);
  k2_1(3) <= out0_66;

  const_expression_19 <= to_unsigned(16#03#, 8);

  out0_75 <= j_j - const_expression_19;

  const_expression_20 <= to_unsigned(16#22#, 8);

  out0_76 <= j_j - const_expression_20;

  const_expression_21 <= to_unsigned(16#02#, 8);

  out0_77 <= j_j - const_expression_21;

  const_expression_22 <= to_unsigned(16#21#, 8);

  out0_78 <= j_j - const_expression_22;

  const_expression_23 <= to_unsigned(16#01#, 8);

  out0_79 <= j_j - const_expression_23;

  const_expression_24 <= to_unsigned(16#20#, 8);

  out0_80 <= j_j - const_expression_24;

  const_expression_25 <= to_unsigned(16#00#, 8);

  out0_81 <= j_j - const_expression_25;

  key_signal1_unsigned <= unsigned(key_signal1);

  Delay5_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal1 <= key_signal1_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_1_process;


  key_signal2_unsigned <= unsigned(key_signal2);

  Delay5_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal2 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal2 <= key_signal2_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_2_process;


  key_signal3_unsigned <= unsigned(key_signal3);

  Delay5_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal3 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal3 <= key_signal3_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_3_process;


  key_signal4_unsigned <= unsigned(key_signal4);

  Delay5_4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal4 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal4 <= key_signal4_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_4_process;


  key_signal5_unsigned <= unsigned(key_signal5);

  Delay5_5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal5 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal5 <= key_signal5_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_5_process;


  key_signal6_unsigned <= unsigned(key_signal6);

  Delay5_6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal6 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal6 <= key_signal6_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_6_process;


  key_signal7_unsigned <= unsigned(key_signal7);

  Delay5_7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal7 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal7 <= key_signal7_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_7_process;


  key_signal8_unsigned <= unsigned(key_signal8);

  Delay5_8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal8 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal8 <= key_signal8_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_8_process;


  key_signal9_unsigned <= unsigned(key_signal9);

  Delay5_9_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal9 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal9 <= key_signal9_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_9_process;


  key_signal10_unsigned <= unsigned(key_signal10);

  Delay5_10_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal10 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal10 <= key_signal10_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_10_process;


  key_signal11_unsigned <= unsigned(key_signal11);

  Delay5_11_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal11 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal11 <= key_signal11_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_11_process;


  key_signal12_unsigned <= unsigned(key_signal12);

  Delay5_12_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal12 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal12 <= key_signal12_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_12_process;


  key_signal13_unsigned <= unsigned(key_signal13);

  Delay5_13_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal13 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal13 <= key_signal13_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_13_process;


  key_signal14_unsigned <= unsigned(key_signal14);

  Delay5_14_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal14 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal14 <= key_signal14_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_14_process;


  key_signal15_unsigned <= unsigned(key_signal15);

  Delay5_15_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal15 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal15 <= key_signal15_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_15_process;


  key_signal16_unsigned <= unsigned(key_signal16);

  Delay5_16_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal16 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal16 <= key_signal16_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_16_process;


  key_signal17_unsigned <= unsigned(key_signal17);

  Delay5_17_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal17 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal17 <= key_signal17_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_17_process;


  key_signal18_unsigned <= unsigned(key_signal18);

  Delay5_18_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal18 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal18 <= key_signal18_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_18_process;


  key_signal19_unsigned <= unsigned(key_signal19);

  Delay5_19_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal19 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal19 <= key_signal19_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_19_process;


  key_signal20_unsigned <= unsigned(key_signal20);

  Delay5_20_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal20 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal20 <= key_signal20_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_20_process;


  key_signal21_unsigned <= unsigned(key_signal21);

  Delay5_21_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal21 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal21 <= key_signal21_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_21_process;


  key_signal22_unsigned <= unsigned(key_signal22);

  Delay5_22_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal22 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal22 <= key_signal22_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_22_process;


  key_signal23_unsigned <= unsigned(key_signal23);

  Delay5_23_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal23 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal23 <= key_signal23_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_23_process;


  key_signal24_unsigned <= unsigned(key_signal24);

  Delay5_24_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal24 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal24 <= key_signal24_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_24_process;


  key_signal25_unsigned <= unsigned(key_signal25);

  Delay5_25_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal25 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal25 <= key_signal25_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_25_process;


  key_signal26_unsigned <= unsigned(key_signal26);

  Delay5_26_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal26 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal26 <= key_signal26_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_26_process;


  key_signal27_unsigned <= unsigned(key_signal27);

  Delay5_27_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal27 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal27 <= key_signal27_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_27_process;


  key_signal28_unsigned <= unsigned(key_signal28);

  Delay5_28_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal28 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal28 <= key_signal28_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_28_process;


  key_signal29_unsigned <= unsigned(key_signal29);

  Delay5_29_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal29 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal29 <= key_signal29_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_29_process;


  key_signal30_unsigned <= unsigned(key_signal30);

  Delay5_30_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal30 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal30 <= key_signal30_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_30_process;


  key_signal31_unsigned <= unsigned(key_signal31);

  Delay5_31_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal31 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal31 <= key_signal31_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_31_process;


  key_signal32_unsigned <= unsigned(key_signal32);

  Delay5_32_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal32 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal32 <= key_signal32_unsigned;
      END IF;
    END IF;
  END PROCESS Delay5_32_process;


  Delay5_out1_to_vector(0) <= signal1;
  Delay5_out1_to_vector(1) <= signal2;
  Delay5_out1_to_vector(2) <= signal3;
  Delay5_out1_to_vector(3) <= signal4;
  Delay5_out1_to_vector(4) <= signal5;
  Delay5_out1_to_vector(5) <= signal6;
  Delay5_out1_to_vector(6) <= signal7;
  Delay5_out1_to_vector(7) <= signal8;
  Delay5_out1_to_vector(8) <= signal9;
  Delay5_out1_to_vector(9) <= signal10;
  Delay5_out1_to_vector(10) <= signal11;
  Delay5_out1_to_vector(11) <= signal12;
  Delay5_out1_to_vector(12) <= signal13;
  Delay5_out1_to_vector(13) <= signal14;
  Delay5_out1_to_vector(14) <= signal15;
  Delay5_out1_to_vector(15) <= signal16;
  Delay5_out1_to_vector(16) <= signal17;
  Delay5_out1_to_vector(17) <= signal18;
  Delay5_out1_to_vector(18) <= signal19;
  Delay5_out1_to_vector(19) <= signal20;
  Delay5_out1_to_vector(20) <= signal21;
  Delay5_out1_to_vector(21) <= signal22;
  Delay5_out1_to_vector(22) <= signal23;
  Delay5_out1_to_vector(23) <= signal24;
  Delay5_out1_to_vector(24) <= signal25;
  Delay5_out1_to_vector(25) <= signal26;
  Delay5_out1_to_vector(26) <= signal27;
  Delay5_out1_to_vector(27) <= signal28;
  Delay5_out1_to_vector(28) <= signal29;
  Delay5_out1_to_vector(29) <= signal30;
  Delay5_out1_to_vector(30) <= signal31;
  Delay5_out1_to_vector(31) <= signal32;

  expandedKey_1(0) <= Delay5_out1_to_vector(0);
  expandedKey_1(1) <= Delay5_out1_to_vector(1);
  expandedKey_1(2) <= Delay5_out1_to_vector(2);
  expandedKey_1(3) <= Delay5_out1_to_vector(3);
  expandedKey_1(4) <= Delay5_out1_to_vector(4);
  expandedKey_1(5) <= Delay5_out1_to_vector(5);
  expandedKey_1(6) <= Delay5_out1_to_vector(6);
  expandedKey_1(7) <= Delay5_out1_to_vector(7);
  expandedKey_1(8) <= Delay5_out1_to_vector(8);
  expandedKey_1(9) <= Delay5_out1_to_vector(9);
  expandedKey_1(10) <= Delay5_out1_to_vector(10);
  expandedKey_1(11) <= Delay5_out1_to_vector(11);
  expandedKey_1(12) <= Delay5_out1_to_vector(12);
  expandedKey_1(13) <= Delay5_out1_to_vector(13);
  expandedKey_1(14) <= Delay5_out1_to_vector(14);
  expandedKey_1(15) <= Delay5_out1_to_vector(15);
  expandedKey_1(16) <= Delay5_out1_to_vector(16);
  expandedKey_1(17) <= Delay5_out1_to_vector(17);
  expandedKey_1(18) <= Delay5_out1_to_vector(18);
  expandedKey_1(19) <= Delay5_out1_to_vector(19);
  expandedKey_1(20) <= Delay5_out1_to_vector(20);
  expandedKey_1(21) <= Delay5_out1_to_vector(21);
  expandedKey_1(22) <= Delay5_out1_to_vector(22);
  expandedKey_1(23) <= Delay5_out1_to_vector(23);
  expandedKey_1(24) <= Delay5_out1_to_vector(24);
  expandedKey_1(25) <= Delay5_out1_to_vector(25);
  expandedKey_1(26) <= Delay5_out1_to_vector(26);
  expandedKey_1(27) <= Delay5_out1_to_vector(27);
  expandedKey_1(28) <= Delay5_out1_to_vector(28);
  expandedKey_1(29) <= Delay5_out1_to_vector(29);
  expandedKey_1(30) <= Delay5_out1_to_vector(30);
  expandedKey_1(31) <= Delay5_out1_to_vector(31);
  expandedKey_1(32) <= expandedKey(32);
  expandedKey_1(33) <= expandedKey(33);
  expandedKey_1(34) <= expandedKey(34);
  expandedKey_1(35) <= expandedKey(35);
  expandedKey_1(36) <= expandedKey(36);
  expandedKey_1(37) <= expandedKey(37);
  expandedKey_1(38) <= expandedKey(38);
  expandedKey_1(39) <= expandedKey(39);
  expandedKey_1(40) <= expandedKey(40);
  expandedKey_1(41) <= expandedKey(41);
  expandedKey_1(42) <= expandedKey(42);
  expandedKey_1(43) <= expandedKey(43);
  expandedKey_1(44) <= expandedKey(44);
  expandedKey_1(45) <= expandedKey(45);
  expandedKey_1(46) <= expandedKey(46);
  expandedKey_1(47) <= expandedKey(47);
  expandedKey_1(48) <= expandedKey(48);
  expandedKey_1(49) <= expandedKey(49);
  expandedKey_1(50) <= expandedKey(50);
  expandedKey_1(51) <= expandedKey(51);
  expandedKey_1(52) <= expandedKey(52);
  expandedKey_1(53) <= expandedKey(53);
  expandedKey_1(54) <= expandedKey(54);
  expandedKey_1(55) <= expandedKey(55);
  expandedKey_1(56) <= expandedKey(56);
  expandedKey_1(57) <= expandedKey(57);
  expandedKey_1(58) <= expandedKey(58);
  expandedKey_1(59) <= expandedKey(59);
  expandedKey_1(60) <= expandedKey(60);
  expandedKey_1(61) <= expandedKey(61);
  expandedKey_1(62) <= expandedKey(62);
  expandedKey_1(63) <= expandedKey(63);
  expandedKey_1(64) <= expandedKey(64);
  expandedKey_1(65) <= expandedKey(65);
  expandedKey_1(66) <= expandedKey(66);
  expandedKey_1(67) <= expandedKey(67);
  expandedKey_1(68) <= expandedKey(68);
  expandedKey_1(69) <= expandedKey(69);
  expandedKey_1(70) <= expandedKey(70);
  expandedKey_1(71) <= expandedKey(71);
  expandedKey_1(72) <= expandedKey(72);
  expandedKey_1(73) <= expandedKey(73);
  expandedKey_1(74) <= expandedKey(74);
  expandedKey_1(75) <= expandedKey(75);
  expandedKey_1(76) <= expandedKey(76);
  expandedKey_1(77) <= expandedKey(77);
  expandedKey_1(78) <= expandedKey(78);
  expandedKey_1(79) <= expandedKey(79);
  expandedKey_1(80) <= expandedKey(80);
  expandedKey_1(81) <= expandedKey(81);
  expandedKey_1(82) <= expandedKey(82);
  expandedKey_1(83) <= expandedKey(83);
  expandedKey_1(84) <= expandedKey(84);
  expandedKey_1(85) <= expandedKey(85);
  expandedKey_1(86) <= expandedKey(86);
  expandedKey_1(87) <= expandedKey(87);
  expandedKey_1(88) <= expandedKey(88);
  expandedKey_1(89) <= expandedKey(89);
  expandedKey_1(90) <= expandedKey(90);
  expandedKey_1(91) <= expandedKey(91);
  expandedKey_1(92) <= expandedKey(92);
  expandedKey_1(93) <= expandedKey(93);
  expandedKey_1(94) <= expandedKey(94);
  expandedKey_1(95) <= expandedKey(95);
  expandedKey_1(96) <= expandedKey(96);
  expandedKey_1(97) <= expandedKey(97);
  expandedKey_1(98) <= expandedKey(98);
  expandedKey_1(99) <= expandedKey(99);
  expandedKey_1(100) <= expandedKey(100);
  expandedKey_1(101) <= expandedKey(101);
  expandedKey_1(102) <= expandedKey(102);
  expandedKey_1(103) <= expandedKey(103);
  expandedKey_1(104) <= expandedKey(104);
  expandedKey_1(105) <= expandedKey(105);
  expandedKey_1(106) <= expandedKey(106);
  expandedKey_1(107) <= expandedKey(107);
  expandedKey_1(108) <= expandedKey(108);
  expandedKey_1(109) <= expandedKey(109);
  expandedKey_1(110) <= expandedKey(110);
  expandedKey_1(111) <= expandedKey(111);
  expandedKey_1(112) <= expandedKey(112);
  expandedKey_1(113) <= expandedKey(113);
  expandedKey_1(114) <= expandedKey(114);
  expandedKey_1(115) <= expandedKey(115);
  expandedKey_1(116) <= expandedKey(116);
  expandedKey_1(117) <= expandedKey(117);
  expandedKey_1(118) <= expandedKey(118);
  expandedKey_1(119) <= expandedKey(119);
  expandedKey_1(120) <= expandedKey(120);
  expandedKey_1(121) <= expandedKey(121);
  expandedKey_1(122) <= expandedKey(122);
  expandedKey_1(123) <= expandedKey(123);
  expandedKey_1(124) <= expandedKey(124);
  expandedKey_1(125) <= expandedKey(125);
  expandedKey_1(126) <= expandedKey(126);
  expandedKey_1(127) <= expandedKey(127);
  expandedKey_1(128) <= expandedKey(128);
  expandedKey_1(129) <= expandedKey(129);
  expandedKey_1(130) <= expandedKey(130);
  expandedKey_1(131) <= expandedKey(131);
  expandedKey_1(132) <= expandedKey(132);
  expandedKey_1(133) <= expandedKey(133);
  expandedKey_1(134) <= expandedKey(134);
  expandedKey_1(135) <= expandedKey(135);
  expandedKey_1(136) <= expandedKey(136);
  expandedKey_1(137) <= expandedKey(137);
  expandedKey_1(138) <= expandedKey(138);
  expandedKey_1(139) <= expandedKey(139);
  expandedKey_1(140) <= expandedKey(140);
  expandedKey_1(141) <= expandedKey(141);
  expandedKey_1(142) <= expandedKey(142);
  expandedKey_1(143) <= expandedKey(143);
  expandedKey_1(144) <= expandedKey(144);
  expandedKey_1(145) <= expandedKey(145);
  expandedKey_1(146) <= expandedKey(146);
  expandedKey_1(147) <= expandedKey(147);
  expandedKey_1(148) <= expandedKey(148);
  expandedKey_1(149) <= expandedKey(149);
  expandedKey_1(150) <= expandedKey(150);
  expandedKey_1(151) <= expandedKey(151);
  expandedKey_1(152) <= expandedKey(152);
  expandedKey_1(153) <= expandedKey(153);
  expandedKey_1(154) <= expandedKey(154);
  expandedKey_1(155) <= expandedKey(155);
  expandedKey_1(156) <= expandedKey(156);
  expandedKey_1(157) <= expandedKey(157);
  expandedKey_1(158) <= expandedKey(158);
  expandedKey_1(159) <= expandedKey(159);
  expandedKey_1(160) <= expandedKey(160);
  expandedKey_1(161) <= expandedKey(161);
  expandedKey_1(162) <= expandedKey(162);
  expandedKey_1(163) <= expandedKey(163);
  expandedKey_1(164) <= expandedKey(164);
  expandedKey_1(165) <= expandedKey(165);
  expandedKey_1(166) <= expandedKey(166);
  expandedKey_1(167) <= expandedKey(167);
  expandedKey_1(168) <= expandedKey(168);
  expandedKey_1(169) <= expandedKey(169);
  expandedKey_1(170) <= expandedKey(170);
  expandedKey_1(171) <= expandedKey(171);
  expandedKey_1(172) <= expandedKey(172);
  expandedKey_1(173) <= expandedKey(173);
  expandedKey_1(174) <= expandedKey(174);
  expandedKey_1(175) <= expandedKey(175);
  expandedKey_1(176) <= expandedKey(176);
  expandedKey_1(177) <= expandedKey(177);
  expandedKey_1(178) <= expandedKey(178);
  expandedKey_1(179) <= expandedKey(179);
  expandedKey_1(180) <= expandedKey(180);
  expandedKey_1(181) <= expandedKey(181);
  expandedKey_1(182) <= expandedKey(182);
  expandedKey_1(183) <= expandedKey(183);
  expandedKey_1(184) <= expandedKey(184);
  expandedKey_1(185) <= expandedKey(185);
  expandedKey_1(186) <= expandedKey(186);
  expandedKey_1(187) <= expandedKey(187);
  expandedKey_1(188) <= expandedKey(188);
  expandedKey_1(189) <= expandedKey(189);
  expandedKey_1(190) <= expandedKey(190);
  expandedKey_1(191) <= expandedKey(191);
  expandedKey_1(192) <= expandedKey(192);
  expandedKey_1(193) <= expandedKey(193);
  expandedKey_1(194) <= expandedKey(194);
  expandedKey_1(195) <= expandedKey(195);
  expandedKey_1(196) <= expandedKey(196);
  expandedKey_1(197) <= expandedKey(197);
  expandedKey_1(198) <= expandedKey(198);
  expandedKey_1(199) <= expandedKey(199);
  expandedKey_1(200) <= expandedKey(200);
  expandedKey_1(201) <= expandedKey(201);
  expandedKey_1(202) <= expandedKey(202);
  expandedKey_1(203) <= expandedKey(203);
  expandedKey_1(204) <= expandedKey(204);
  expandedKey_1(205) <= expandedKey(205);
  expandedKey_1(206) <= expandedKey(206);
  expandedKey_1(207) <= expandedKey(207);
  expandedKey_1(208) <= expandedKey(208);
  expandedKey_1(209) <= expandedKey(209);
  expandedKey_1(210) <= expandedKey(210);
  expandedKey_1(211) <= expandedKey(211);
  expandedKey_1(212) <= expandedKey(212);
  expandedKey_1(213) <= expandedKey(213);
  expandedKey_1(214) <= expandedKey(214);
  expandedKey_1(215) <= expandedKey(215);
  expandedKey_1(216) <= expandedKey(216);
  expandedKey_1(217) <= expandedKey(217);
  expandedKey_1(218) <= expandedKey(218);
  expandedKey_1(219) <= expandedKey(219);
  expandedKey_1(220) <= expandedKey(220);
  expandedKey_1(221) <= expandedKey(221);
  expandedKey_1(222) <= expandedKey(222);
  expandedKey_1(223) <= expandedKey(223);
  expandedKey_1(224) <= expandedKey(224);
  expandedKey_1(225) <= expandedKey(225);
  expandedKey_1(226) <= expandedKey(226);
  expandedKey_1(227) <= expandedKey(227);
  expandedKey_1(228) <= expandedKey(228);
  expandedKey_1(229) <= expandedKey(229);
  expandedKey_1(230) <= expandedKey(230);
  expandedKey_1(231) <= expandedKey(231);
  expandedKey_1(232) <= expandedKey(232);
  expandedKey_1(233) <= expandedKey(233);
  expandedKey_1(234) <= expandedKey(234);
  expandedKey_1(235) <= expandedKey(235);
  expandedKey_1(236) <= expandedKey(236);
  expandedKey_1(237) <= expandedKey(237);
  expandedKey_1(238) <= expandedKey(238);
  expandedKey_1(239) <= expandedKey(239);

  temp_key_3 <= temp_key(3);

  
  out0_82 <= expandedKey_2(0) WHEN out0_80 = to_unsigned(16#01#, 8) ELSE
      expandedKey_2(1) WHEN out0_80 = to_unsigned(16#02#, 8) ELSE
      expandedKey_2(2) WHEN out0_80 = to_unsigned(16#03#, 8) ELSE
      expandedKey_2(3) WHEN out0_80 = to_unsigned(16#04#, 8) ELSE
      expandedKey_2(4) WHEN out0_80 = to_unsigned(16#05#, 8) ELSE
      expandedKey_2(5) WHEN out0_80 = to_unsigned(16#06#, 8) ELSE
      expandedKey_2(6) WHEN out0_80 = to_unsigned(16#07#, 8) ELSE
      expandedKey_2(7) WHEN out0_80 = to_unsigned(16#08#, 8) ELSE
      expandedKey_2(8) WHEN out0_80 = to_unsigned(16#09#, 8) ELSE
      expandedKey_2(9) WHEN out0_80 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_2(10) WHEN out0_80 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_2(11) WHEN out0_80 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_2(12) WHEN out0_80 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_2(13) WHEN out0_80 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_2(14) WHEN out0_80 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_2(15) WHEN out0_80 = to_unsigned(16#10#, 8) ELSE
      expandedKey_2(16) WHEN out0_80 = to_unsigned(16#11#, 8) ELSE
      expandedKey_2(17) WHEN out0_80 = to_unsigned(16#12#, 8) ELSE
      expandedKey_2(18) WHEN out0_80 = to_unsigned(16#13#, 8) ELSE
      expandedKey_2(19) WHEN out0_80 = to_unsigned(16#14#, 8) ELSE
      expandedKey_2(20) WHEN out0_80 = to_unsigned(16#15#, 8) ELSE
      expandedKey_2(21) WHEN out0_80 = to_unsigned(16#16#, 8) ELSE
      expandedKey_2(22) WHEN out0_80 = to_unsigned(16#17#, 8) ELSE
      expandedKey_2(23) WHEN out0_80 = to_unsigned(16#18#, 8) ELSE
      expandedKey_2(24) WHEN out0_80 = to_unsigned(16#19#, 8) ELSE
      expandedKey_2(25) WHEN out0_80 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_2(26) WHEN out0_80 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_2(27) WHEN out0_80 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_2(28) WHEN out0_80 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_2(29) WHEN out0_80 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_2(30) WHEN out0_80 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_2(31) WHEN out0_80 = to_unsigned(16#20#, 8) ELSE
      expandedKey_2(32) WHEN out0_80 = to_unsigned(16#21#, 8) ELSE
      expandedKey_2(33) WHEN out0_80 = to_unsigned(16#22#, 8) ELSE
      expandedKey_2(34) WHEN out0_80 = to_unsigned(16#23#, 8) ELSE
      expandedKey_2(35) WHEN out0_80 = to_unsigned(16#24#, 8) ELSE
      expandedKey_2(36) WHEN out0_80 = to_unsigned(16#25#, 8) ELSE
      expandedKey_2(37) WHEN out0_80 = to_unsigned(16#26#, 8) ELSE
      expandedKey_2(38) WHEN out0_80 = to_unsigned(16#27#, 8) ELSE
      expandedKey_2(39) WHEN out0_80 = to_unsigned(16#28#, 8) ELSE
      expandedKey_2(40) WHEN out0_80 = to_unsigned(16#29#, 8) ELSE
      expandedKey_2(41) WHEN out0_80 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_2(42) WHEN out0_80 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_2(43) WHEN out0_80 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_2(44) WHEN out0_80 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_2(45) WHEN out0_80 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_2(46) WHEN out0_80 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_2(47) WHEN out0_80 = to_unsigned(16#30#, 8) ELSE
      expandedKey_2(48) WHEN out0_80 = to_unsigned(16#31#, 8) ELSE
      expandedKey_2(49) WHEN out0_80 = to_unsigned(16#32#, 8) ELSE
      expandedKey_2(50) WHEN out0_80 = to_unsigned(16#33#, 8) ELSE
      expandedKey_2(51) WHEN out0_80 = to_unsigned(16#34#, 8) ELSE
      expandedKey_2(52) WHEN out0_80 = to_unsigned(16#35#, 8) ELSE
      expandedKey_2(53) WHEN out0_80 = to_unsigned(16#36#, 8) ELSE
      expandedKey_2(54) WHEN out0_80 = to_unsigned(16#37#, 8) ELSE
      expandedKey_2(55) WHEN out0_80 = to_unsigned(16#38#, 8) ELSE
      expandedKey_2(56) WHEN out0_80 = to_unsigned(16#39#, 8) ELSE
      expandedKey_2(57) WHEN out0_80 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_2(58) WHEN out0_80 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_2(59) WHEN out0_80 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_2(60) WHEN out0_80 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_2(61) WHEN out0_80 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_2(62) WHEN out0_80 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_2(63) WHEN out0_80 = to_unsigned(16#40#, 8) ELSE
      expandedKey_2(64) WHEN out0_80 = to_unsigned(16#41#, 8) ELSE
      expandedKey_2(65) WHEN out0_80 = to_unsigned(16#42#, 8) ELSE
      expandedKey_2(66) WHEN out0_80 = to_unsigned(16#43#, 8) ELSE
      expandedKey_2(67) WHEN out0_80 = to_unsigned(16#44#, 8) ELSE
      expandedKey_2(68) WHEN out0_80 = to_unsigned(16#45#, 8) ELSE
      expandedKey_2(69) WHEN out0_80 = to_unsigned(16#46#, 8) ELSE
      expandedKey_2(70) WHEN out0_80 = to_unsigned(16#47#, 8) ELSE
      expandedKey_2(71) WHEN out0_80 = to_unsigned(16#48#, 8) ELSE
      expandedKey_2(72) WHEN out0_80 = to_unsigned(16#49#, 8) ELSE
      expandedKey_2(73) WHEN out0_80 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_2(74) WHEN out0_80 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_2(75) WHEN out0_80 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_2(76) WHEN out0_80 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_2(77) WHEN out0_80 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_2(78) WHEN out0_80 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_2(79) WHEN out0_80 = to_unsigned(16#50#, 8) ELSE
      expandedKey_2(80) WHEN out0_80 = to_unsigned(16#51#, 8) ELSE
      expandedKey_2(81) WHEN out0_80 = to_unsigned(16#52#, 8) ELSE
      expandedKey_2(82) WHEN out0_80 = to_unsigned(16#53#, 8) ELSE
      expandedKey_2(83) WHEN out0_80 = to_unsigned(16#54#, 8) ELSE
      expandedKey_2(84) WHEN out0_80 = to_unsigned(16#55#, 8) ELSE
      expandedKey_2(85) WHEN out0_80 = to_unsigned(16#56#, 8) ELSE
      expandedKey_2(86) WHEN out0_80 = to_unsigned(16#57#, 8) ELSE
      expandedKey_2(87) WHEN out0_80 = to_unsigned(16#58#, 8) ELSE
      expandedKey_2(88) WHEN out0_80 = to_unsigned(16#59#, 8) ELSE
      expandedKey_2(89) WHEN out0_80 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_2(90) WHEN out0_80 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_2(91) WHEN out0_80 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_2(92) WHEN out0_80 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_2(93) WHEN out0_80 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_2(94) WHEN out0_80 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_2(95) WHEN out0_80 = to_unsigned(16#60#, 8) ELSE
      expandedKey_2(96) WHEN out0_80 = to_unsigned(16#61#, 8) ELSE
      expandedKey_2(97) WHEN out0_80 = to_unsigned(16#62#, 8) ELSE
      expandedKey_2(98) WHEN out0_80 = to_unsigned(16#63#, 8) ELSE
      expandedKey_2(99) WHEN out0_80 = to_unsigned(16#64#, 8) ELSE
      expandedKey_2(100) WHEN out0_80 = to_unsigned(16#65#, 8) ELSE
      expandedKey_2(101) WHEN out0_80 = to_unsigned(16#66#, 8) ELSE
      expandedKey_2(102) WHEN out0_80 = to_unsigned(16#67#, 8) ELSE
      expandedKey_2(103) WHEN out0_80 = to_unsigned(16#68#, 8) ELSE
      expandedKey_2(104) WHEN out0_80 = to_unsigned(16#69#, 8) ELSE
      expandedKey_2(105) WHEN out0_80 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_2(106) WHEN out0_80 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_2(107) WHEN out0_80 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_2(108) WHEN out0_80 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_2(109) WHEN out0_80 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_2(110) WHEN out0_80 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_2(111) WHEN out0_80 = to_unsigned(16#70#, 8) ELSE
      expandedKey_2(112) WHEN out0_80 = to_unsigned(16#71#, 8) ELSE
      expandedKey_2(113) WHEN out0_80 = to_unsigned(16#72#, 8) ELSE
      expandedKey_2(114) WHEN out0_80 = to_unsigned(16#73#, 8) ELSE
      expandedKey_2(115) WHEN out0_80 = to_unsigned(16#74#, 8) ELSE
      expandedKey_2(116) WHEN out0_80 = to_unsigned(16#75#, 8) ELSE
      expandedKey_2(117) WHEN out0_80 = to_unsigned(16#76#, 8) ELSE
      expandedKey_2(118) WHEN out0_80 = to_unsigned(16#77#, 8) ELSE
      expandedKey_2(119) WHEN out0_80 = to_unsigned(16#78#, 8) ELSE
      expandedKey_2(120) WHEN out0_80 = to_unsigned(16#79#, 8) ELSE
      expandedKey_2(121) WHEN out0_80 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_2(122) WHEN out0_80 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_2(123) WHEN out0_80 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_2(124) WHEN out0_80 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_2(125) WHEN out0_80 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_2(126) WHEN out0_80 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_2(127) WHEN out0_80 = to_unsigned(16#80#, 8) ELSE
      expandedKey_2(128) WHEN out0_80 = to_unsigned(16#81#, 8) ELSE
      expandedKey_2(129) WHEN out0_80 = to_unsigned(16#82#, 8) ELSE
      expandedKey_2(130) WHEN out0_80 = to_unsigned(16#83#, 8) ELSE
      expandedKey_2(131) WHEN out0_80 = to_unsigned(16#84#, 8) ELSE
      expandedKey_2(132) WHEN out0_80 = to_unsigned(16#85#, 8) ELSE
      expandedKey_2(133) WHEN out0_80 = to_unsigned(16#86#, 8) ELSE
      expandedKey_2(134) WHEN out0_80 = to_unsigned(16#87#, 8) ELSE
      expandedKey_2(135) WHEN out0_80 = to_unsigned(16#88#, 8) ELSE
      expandedKey_2(136) WHEN out0_80 = to_unsigned(16#89#, 8) ELSE
      expandedKey_2(137) WHEN out0_80 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_2(138) WHEN out0_80 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_2(139) WHEN out0_80 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_2(140) WHEN out0_80 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_2(141) WHEN out0_80 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_2(142) WHEN out0_80 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_2(143) WHEN out0_80 = to_unsigned(16#90#, 8) ELSE
      expandedKey_2(144) WHEN out0_80 = to_unsigned(16#91#, 8) ELSE
      expandedKey_2(145) WHEN out0_80 = to_unsigned(16#92#, 8) ELSE
      expandedKey_2(146) WHEN out0_80 = to_unsigned(16#93#, 8) ELSE
      expandedKey_2(147) WHEN out0_80 = to_unsigned(16#94#, 8) ELSE
      expandedKey_2(148) WHEN out0_80 = to_unsigned(16#95#, 8) ELSE
      expandedKey_2(149) WHEN out0_80 = to_unsigned(16#96#, 8) ELSE
      expandedKey_2(150) WHEN out0_80 = to_unsigned(16#97#, 8) ELSE
      expandedKey_2(151) WHEN out0_80 = to_unsigned(16#98#, 8) ELSE
      expandedKey_2(152) WHEN out0_80 = to_unsigned(16#99#, 8) ELSE
      expandedKey_2(153) WHEN out0_80 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_2(154) WHEN out0_80 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_2(155) WHEN out0_80 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_2(156) WHEN out0_80 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_2(157) WHEN out0_80 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_2(158) WHEN out0_80 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_2(159) WHEN out0_80 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_2(160) WHEN out0_80 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_2(161) WHEN out0_80 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_2(162) WHEN out0_80 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_2(163) WHEN out0_80 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_2(164) WHEN out0_80 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_2(165) WHEN out0_80 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_2(166) WHEN out0_80 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_2(167) WHEN out0_80 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_2(168) WHEN out0_80 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_2(169) WHEN out0_80 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_2(170) WHEN out0_80 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_2(171) WHEN out0_80 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_2(172) WHEN out0_80 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_2(173) WHEN out0_80 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_2(174) WHEN out0_80 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_2(175) WHEN out0_80 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_2(176) WHEN out0_80 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_2(177) WHEN out0_80 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_2(178) WHEN out0_80 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_2(179) WHEN out0_80 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_2(180) WHEN out0_80 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_2(181) WHEN out0_80 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_2(182) WHEN out0_80 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_2(183) WHEN out0_80 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_2(184) WHEN out0_80 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_2(185) WHEN out0_80 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_2(186) WHEN out0_80 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_2(187) WHEN out0_80 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_2(188) WHEN out0_80 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_2(189) WHEN out0_80 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_2(190) WHEN out0_80 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_2(191) WHEN out0_80 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_2(192) WHEN out0_80 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_2(193) WHEN out0_80 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_2(194) WHEN out0_80 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_2(195) WHEN out0_80 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_2(196) WHEN out0_80 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_2(197) WHEN out0_80 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_2(198) WHEN out0_80 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_2(199) WHEN out0_80 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_2(200) WHEN out0_80 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_2(201) WHEN out0_80 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_2(202) WHEN out0_80 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_2(203) WHEN out0_80 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_2(204) WHEN out0_80 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_2(205) WHEN out0_80 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_2(206) WHEN out0_80 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_2(207) WHEN out0_80 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_2(208) WHEN out0_80 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_2(209) WHEN out0_80 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_2(210) WHEN out0_80 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_2(211) WHEN out0_80 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_2(212) WHEN out0_80 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_2(213) WHEN out0_80 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_2(214) WHEN out0_80 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_2(215) WHEN out0_80 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_2(216) WHEN out0_80 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_2(217) WHEN out0_80 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_2(218) WHEN out0_80 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_2(219) WHEN out0_80 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_2(220) WHEN out0_80 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_2(221) WHEN out0_80 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_2(222) WHEN out0_80 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_2(223) WHEN out0_80 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_2(224) WHEN out0_80 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_2(225) WHEN out0_80 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_2(226) WHEN out0_80 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_2(227) WHEN out0_80 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_2(228) WHEN out0_80 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_2(229) WHEN out0_80 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_2(230) WHEN out0_80 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_2(231) WHEN out0_80 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_2(232) WHEN out0_80 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_2(233) WHEN out0_80 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_2(234) WHEN out0_80 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_2(235) WHEN out0_80 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_2(236) WHEN out0_80 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_2(237) WHEN out0_80 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_2(238) WHEN out0_80 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_2(239);

  out0_83 <= out0_82 XOR temp_key_3;

  temp_key_2 <= temp_key(2);

  
  out0_84 <= expandedKey_3(0) WHEN out0_78 = to_unsigned(16#01#, 8) ELSE
      expandedKey_3(1) WHEN out0_78 = to_unsigned(16#02#, 8) ELSE
      expandedKey_3(2) WHEN out0_78 = to_unsigned(16#03#, 8) ELSE
      expandedKey_3(3) WHEN out0_78 = to_unsigned(16#04#, 8) ELSE
      expandedKey_3(4) WHEN out0_78 = to_unsigned(16#05#, 8) ELSE
      expandedKey_3(5) WHEN out0_78 = to_unsigned(16#06#, 8) ELSE
      expandedKey_3(6) WHEN out0_78 = to_unsigned(16#07#, 8) ELSE
      expandedKey_3(7) WHEN out0_78 = to_unsigned(16#08#, 8) ELSE
      expandedKey_3(8) WHEN out0_78 = to_unsigned(16#09#, 8) ELSE
      expandedKey_3(9) WHEN out0_78 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_3(10) WHEN out0_78 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_3(11) WHEN out0_78 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_3(12) WHEN out0_78 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_3(13) WHEN out0_78 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_3(14) WHEN out0_78 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_3(15) WHEN out0_78 = to_unsigned(16#10#, 8) ELSE
      expandedKey_3(16) WHEN out0_78 = to_unsigned(16#11#, 8) ELSE
      expandedKey_3(17) WHEN out0_78 = to_unsigned(16#12#, 8) ELSE
      expandedKey_3(18) WHEN out0_78 = to_unsigned(16#13#, 8) ELSE
      expandedKey_3(19) WHEN out0_78 = to_unsigned(16#14#, 8) ELSE
      expandedKey_3(20) WHEN out0_78 = to_unsigned(16#15#, 8) ELSE
      expandedKey_3(21) WHEN out0_78 = to_unsigned(16#16#, 8) ELSE
      expandedKey_3(22) WHEN out0_78 = to_unsigned(16#17#, 8) ELSE
      expandedKey_3(23) WHEN out0_78 = to_unsigned(16#18#, 8) ELSE
      expandedKey_3(24) WHEN out0_78 = to_unsigned(16#19#, 8) ELSE
      expandedKey_3(25) WHEN out0_78 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_3(26) WHEN out0_78 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_3(27) WHEN out0_78 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_3(28) WHEN out0_78 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_3(29) WHEN out0_78 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_3(30) WHEN out0_78 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_3(31) WHEN out0_78 = to_unsigned(16#20#, 8) ELSE
      expandedKey_3(32) WHEN out0_78 = to_unsigned(16#21#, 8) ELSE
      expandedKey_3(33) WHEN out0_78 = to_unsigned(16#22#, 8) ELSE
      expandedKey_3(34) WHEN out0_78 = to_unsigned(16#23#, 8) ELSE
      expandedKey_3(35) WHEN out0_78 = to_unsigned(16#24#, 8) ELSE
      expandedKey_3(36) WHEN out0_78 = to_unsigned(16#25#, 8) ELSE
      expandedKey_3(37) WHEN out0_78 = to_unsigned(16#26#, 8) ELSE
      expandedKey_3(38) WHEN out0_78 = to_unsigned(16#27#, 8) ELSE
      expandedKey_3(39) WHEN out0_78 = to_unsigned(16#28#, 8) ELSE
      expandedKey_3(40) WHEN out0_78 = to_unsigned(16#29#, 8) ELSE
      expandedKey_3(41) WHEN out0_78 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_3(42) WHEN out0_78 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_3(43) WHEN out0_78 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_3(44) WHEN out0_78 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_3(45) WHEN out0_78 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_3(46) WHEN out0_78 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_3(47) WHEN out0_78 = to_unsigned(16#30#, 8) ELSE
      expandedKey_3(48) WHEN out0_78 = to_unsigned(16#31#, 8) ELSE
      expandedKey_3(49) WHEN out0_78 = to_unsigned(16#32#, 8) ELSE
      expandedKey_3(50) WHEN out0_78 = to_unsigned(16#33#, 8) ELSE
      expandedKey_3(51) WHEN out0_78 = to_unsigned(16#34#, 8) ELSE
      expandedKey_3(52) WHEN out0_78 = to_unsigned(16#35#, 8) ELSE
      expandedKey_3(53) WHEN out0_78 = to_unsigned(16#36#, 8) ELSE
      expandedKey_3(54) WHEN out0_78 = to_unsigned(16#37#, 8) ELSE
      expandedKey_3(55) WHEN out0_78 = to_unsigned(16#38#, 8) ELSE
      expandedKey_3(56) WHEN out0_78 = to_unsigned(16#39#, 8) ELSE
      expandedKey_3(57) WHEN out0_78 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_3(58) WHEN out0_78 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_3(59) WHEN out0_78 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_3(60) WHEN out0_78 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_3(61) WHEN out0_78 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_3(62) WHEN out0_78 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_3(63) WHEN out0_78 = to_unsigned(16#40#, 8) ELSE
      expandedKey_3(64) WHEN out0_78 = to_unsigned(16#41#, 8) ELSE
      expandedKey_3(65) WHEN out0_78 = to_unsigned(16#42#, 8) ELSE
      expandedKey_3(66) WHEN out0_78 = to_unsigned(16#43#, 8) ELSE
      expandedKey_3(67) WHEN out0_78 = to_unsigned(16#44#, 8) ELSE
      expandedKey_3(68) WHEN out0_78 = to_unsigned(16#45#, 8) ELSE
      expandedKey_3(69) WHEN out0_78 = to_unsigned(16#46#, 8) ELSE
      expandedKey_3(70) WHEN out0_78 = to_unsigned(16#47#, 8) ELSE
      expandedKey_3(71) WHEN out0_78 = to_unsigned(16#48#, 8) ELSE
      expandedKey_3(72) WHEN out0_78 = to_unsigned(16#49#, 8) ELSE
      expandedKey_3(73) WHEN out0_78 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_3(74) WHEN out0_78 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_3(75) WHEN out0_78 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_3(76) WHEN out0_78 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_3(77) WHEN out0_78 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_3(78) WHEN out0_78 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_3(79) WHEN out0_78 = to_unsigned(16#50#, 8) ELSE
      expandedKey_3(80) WHEN out0_78 = to_unsigned(16#51#, 8) ELSE
      expandedKey_3(81) WHEN out0_78 = to_unsigned(16#52#, 8) ELSE
      expandedKey_3(82) WHEN out0_78 = to_unsigned(16#53#, 8) ELSE
      expandedKey_3(83) WHEN out0_78 = to_unsigned(16#54#, 8) ELSE
      expandedKey_3(84) WHEN out0_78 = to_unsigned(16#55#, 8) ELSE
      expandedKey_3(85) WHEN out0_78 = to_unsigned(16#56#, 8) ELSE
      expandedKey_3(86) WHEN out0_78 = to_unsigned(16#57#, 8) ELSE
      expandedKey_3(87) WHEN out0_78 = to_unsigned(16#58#, 8) ELSE
      expandedKey_3(88) WHEN out0_78 = to_unsigned(16#59#, 8) ELSE
      expandedKey_3(89) WHEN out0_78 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_3(90) WHEN out0_78 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_3(91) WHEN out0_78 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_3(92) WHEN out0_78 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_3(93) WHEN out0_78 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_3(94) WHEN out0_78 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_3(95) WHEN out0_78 = to_unsigned(16#60#, 8) ELSE
      expandedKey_3(96) WHEN out0_78 = to_unsigned(16#61#, 8) ELSE
      expandedKey_3(97) WHEN out0_78 = to_unsigned(16#62#, 8) ELSE
      expandedKey_3(98) WHEN out0_78 = to_unsigned(16#63#, 8) ELSE
      expandedKey_3(99) WHEN out0_78 = to_unsigned(16#64#, 8) ELSE
      expandedKey_3(100) WHEN out0_78 = to_unsigned(16#65#, 8) ELSE
      expandedKey_3(101) WHEN out0_78 = to_unsigned(16#66#, 8) ELSE
      expandedKey_3(102) WHEN out0_78 = to_unsigned(16#67#, 8) ELSE
      expandedKey_3(103) WHEN out0_78 = to_unsigned(16#68#, 8) ELSE
      expandedKey_3(104) WHEN out0_78 = to_unsigned(16#69#, 8) ELSE
      expandedKey_3(105) WHEN out0_78 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_3(106) WHEN out0_78 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_3(107) WHEN out0_78 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_3(108) WHEN out0_78 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_3(109) WHEN out0_78 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_3(110) WHEN out0_78 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_3(111) WHEN out0_78 = to_unsigned(16#70#, 8) ELSE
      expandedKey_3(112) WHEN out0_78 = to_unsigned(16#71#, 8) ELSE
      expandedKey_3(113) WHEN out0_78 = to_unsigned(16#72#, 8) ELSE
      expandedKey_3(114) WHEN out0_78 = to_unsigned(16#73#, 8) ELSE
      expandedKey_3(115) WHEN out0_78 = to_unsigned(16#74#, 8) ELSE
      expandedKey_3(116) WHEN out0_78 = to_unsigned(16#75#, 8) ELSE
      expandedKey_3(117) WHEN out0_78 = to_unsigned(16#76#, 8) ELSE
      expandedKey_3(118) WHEN out0_78 = to_unsigned(16#77#, 8) ELSE
      expandedKey_3(119) WHEN out0_78 = to_unsigned(16#78#, 8) ELSE
      expandedKey_3(120) WHEN out0_78 = to_unsigned(16#79#, 8) ELSE
      expandedKey_3(121) WHEN out0_78 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_3(122) WHEN out0_78 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_3(123) WHEN out0_78 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_3(124) WHEN out0_78 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_3(125) WHEN out0_78 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_3(126) WHEN out0_78 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_3(127) WHEN out0_78 = to_unsigned(16#80#, 8) ELSE
      expandedKey_3(128) WHEN out0_78 = to_unsigned(16#81#, 8) ELSE
      expandedKey_3(129) WHEN out0_78 = to_unsigned(16#82#, 8) ELSE
      expandedKey_3(130) WHEN out0_78 = to_unsigned(16#83#, 8) ELSE
      expandedKey_3(131) WHEN out0_78 = to_unsigned(16#84#, 8) ELSE
      expandedKey_3(132) WHEN out0_78 = to_unsigned(16#85#, 8) ELSE
      expandedKey_3(133) WHEN out0_78 = to_unsigned(16#86#, 8) ELSE
      expandedKey_3(134) WHEN out0_78 = to_unsigned(16#87#, 8) ELSE
      expandedKey_3(135) WHEN out0_78 = to_unsigned(16#88#, 8) ELSE
      expandedKey_3(136) WHEN out0_78 = to_unsigned(16#89#, 8) ELSE
      expandedKey_3(137) WHEN out0_78 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_3(138) WHEN out0_78 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_3(139) WHEN out0_78 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_3(140) WHEN out0_78 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_3(141) WHEN out0_78 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_3(142) WHEN out0_78 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_3(143) WHEN out0_78 = to_unsigned(16#90#, 8) ELSE
      expandedKey_3(144) WHEN out0_78 = to_unsigned(16#91#, 8) ELSE
      expandedKey_3(145) WHEN out0_78 = to_unsigned(16#92#, 8) ELSE
      expandedKey_3(146) WHEN out0_78 = to_unsigned(16#93#, 8) ELSE
      expandedKey_3(147) WHEN out0_78 = to_unsigned(16#94#, 8) ELSE
      expandedKey_3(148) WHEN out0_78 = to_unsigned(16#95#, 8) ELSE
      expandedKey_3(149) WHEN out0_78 = to_unsigned(16#96#, 8) ELSE
      expandedKey_3(150) WHEN out0_78 = to_unsigned(16#97#, 8) ELSE
      expandedKey_3(151) WHEN out0_78 = to_unsigned(16#98#, 8) ELSE
      expandedKey_3(152) WHEN out0_78 = to_unsigned(16#99#, 8) ELSE
      expandedKey_3(153) WHEN out0_78 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_3(154) WHEN out0_78 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_3(155) WHEN out0_78 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_3(156) WHEN out0_78 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_3(157) WHEN out0_78 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_3(158) WHEN out0_78 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_3(159) WHEN out0_78 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_3(160) WHEN out0_78 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_3(161) WHEN out0_78 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_3(162) WHEN out0_78 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_3(163) WHEN out0_78 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_3(164) WHEN out0_78 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_3(165) WHEN out0_78 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_3(166) WHEN out0_78 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_3(167) WHEN out0_78 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_3(168) WHEN out0_78 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_3(169) WHEN out0_78 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_3(170) WHEN out0_78 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_3(171) WHEN out0_78 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_3(172) WHEN out0_78 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_3(173) WHEN out0_78 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_3(174) WHEN out0_78 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_3(175) WHEN out0_78 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_3(176) WHEN out0_78 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_3(177) WHEN out0_78 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_3(178) WHEN out0_78 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_3(179) WHEN out0_78 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_3(180) WHEN out0_78 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_3(181) WHEN out0_78 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_3(182) WHEN out0_78 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_3(183) WHEN out0_78 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_3(184) WHEN out0_78 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_3(185) WHEN out0_78 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_3(186) WHEN out0_78 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_3(187) WHEN out0_78 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_3(188) WHEN out0_78 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_3(189) WHEN out0_78 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_3(190) WHEN out0_78 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_3(191) WHEN out0_78 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_3(192) WHEN out0_78 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_3(193) WHEN out0_78 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_3(194) WHEN out0_78 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_3(195) WHEN out0_78 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_3(196) WHEN out0_78 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_3(197) WHEN out0_78 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_3(198) WHEN out0_78 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_3(199) WHEN out0_78 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_3(200) WHEN out0_78 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_3(201) WHEN out0_78 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_3(202) WHEN out0_78 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_3(203) WHEN out0_78 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_3(204) WHEN out0_78 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_3(205) WHEN out0_78 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_3(206) WHEN out0_78 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_3(207) WHEN out0_78 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_3(208) WHEN out0_78 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_3(209) WHEN out0_78 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_3(210) WHEN out0_78 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_3(211) WHEN out0_78 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_3(212) WHEN out0_78 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_3(213) WHEN out0_78 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_3(214) WHEN out0_78 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_3(215) WHEN out0_78 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_3(216) WHEN out0_78 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_3(217) WHEN out0_78 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_3(218) WHEN out0_78 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_3(219) WHEN out0_78 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_3(220) WHEN out0_78 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_3(221) WHEN out0_78 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_3(222) WHEN out0_78 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_3(223) WHEN out0_78 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_3(224) WHEN out0_78 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_3(225) WHEN out0_78 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_3(226) WHEN out0_78 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_3(227) WHEN out0_78 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_3(228) WHEN out0_78 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_3(229) WHEN out0_78 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_3(230) WHEN out0_78 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_3(231) WHEN out0_78 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_3(232) WHEN out0_78 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_3(233) WHEN out0_78 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_3(234) WHEN out0_78 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_3(235) WHEN out0_78 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_3(236) WHEN out0_78 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_3(237) WHEN out0_78 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_3(238) WHEN out0_78 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_3(239);

  out0_85 <= out0_84 XOR temp_key_2;

  temp_key_1 <= temp_key(1);

  
  out0_86 <= expandedKey_4(0) WHEN out0_76 = to_unsigned(16#01#, 8) ELSE
      expandedKey_4(1) WHEN out0_76 = to_unsigned(16#02#, 8) ELSE
      expandedKey_4(2) WHEN out0_76 = to_unsigned(16#03#, 8) ELSE
      expandedKey_4(3) WHEN out0_76 = to_unsigned(16#04#, 8) ELSE
      expandedKey_4(4) WHEN out0_76 = to_unsigned(16#05#, 8) ELSE
      expandedKey_4(5) WHEN out0_76 = to_unsigned(16#06#, 8) ELSE
      expandedKey_4(6) WHEN out0_76 = to_unsigned(16#07#, 8) ELSE
      expandedKey_4(7) WHEN out0_76 = to_unsigned(16#08#, 8) ELSE
      expandedKey_4(8) WHEN out0_76 = to_unsigned(16#09#, 8) ELSE
      expandedKey_4(9) WHEN out0_76 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_4(10) WHEN out0_76 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_4(11) WHEN out0_76 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_4(12) WHEN out0_76 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_4(13) WHEN out0_76 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_4(14) WHEN out0_76 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_4(15) WHEN out0_76 = to_unsigned(16#10#, 8) ELSE
      expandedKey_4(16) WHEN out0_76 = to_unsigned(16#11#, 8) ELSE
      expandedKey_4(17) WHEN out0_76 = to_unsigned(16#12#, 8) ELSE
      expandedKey_4(18) WHEN out0_76 = to_unsigned(16#13#, 8) ELSE
      expandedKey_4(19) WHEN out0_76 = to_unsigned(16#14#, 8) ELSE
      expandedKey_4(20) WHEN out0_76 = to_unsigned(16#15#, 8) ELSE
      expandedKey_4(21) WHEN out0_76 = to_unsigned(16#16#, 8) ELSE
      expandedKey_4(22) WHEN out0_76 = to_unsigned(16#17#, 8) ELSE
      expandedKey_4(23) WHEN out0_76 = to_unsigned(16#18#, 8) ELSE
      expandedKey_4(24) WHEN out0_76 = to_unsigned(16#19#, 8) ELSE
      expandedKey_4(25) WHEN out0_76 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_4(26) WHEN out0_76 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_4(27) WHEN out0_76 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_4(28) WHEN out0_76 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_4(29) WHEN out0_76 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_4(30) WHEN out0_76 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_4(31) WHEN out0_76 = to_unsigned(16#20#, 8) ELSE
      expandedKey_4(32) WHEN out0_76 = to_unsigned(16#21#, 8) ELSE
      expandedKey_4(33) WHEN out0_76 = to_unsigned(16#22#, 8) ELSE
      expandedKey_4(34) WHEN out0_76 = to_unsigned(16#23#, 8) ELSE
      expandedKey_4(35) WHEN out0_76 = to_unsigned(16#24#, 8) ELSE
      expandedKey_4(36) WHEN out0_76 = to_unsigned(16#25#, 8) ELSE
      expandedKey_4(37) WHEN out0_76 = to_unsigned(16#26#, 8) ELSE
      expandedKey_4(38) WHEN out0_76 = to_unsigned(16#27#, 8) ELSE
      expandedKey_4(39) WHEN out0_76 = to_unsigned(16#28#, 8) ELSE
      expandedKey_4(40) WHEN out0_76 = to_unsigned(16#29#, 8) ELSE
      expandedKey_4(41) WHEN out0_76 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_4(42) WHEN out0_76 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_4(43) WHEN out0_76 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_4(44) WHEN out0_76 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_4(45) WHEN out0_76 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_4(46) WHEN out0_76 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_4(47) WHEN out0_76 = to_unsigned(16#30#, 8) ELSE
      expandedKey_4(48) WHEN out0_76 = to_unsigned(16#31#, 8) ELSE
      expandedKey_4(49) WHEN out0_76 = to_unsigned(16#32#, 8) ELSE
      expandedKey_4(50) WHEN out0_76 = to_unsigned(16#33#, 8) ELSE
      expandedKey_4(51) WHEN out0_76 = to_unsigned(16#34#, 8) ELSE
      expandedKey_4(52) WHEN out0_76 = to_unsigned(16#35#, 8) ELSE
      expandedKey_4(53) WHEN out0_76 = to_unsigned(16#36#, 8) ELSE
      expandedKey_4(54) WHEN out0_76 = to_unsigned(16#37#, 8) ELSE
      expandedKey_4(55) WHEN out0_76 = to_unsigned(16#38#, 8) ELSE
      expandedKey_4(56) WHEN out0_76 = to_unsigned(16#39#, 8) ELSE
      expandedKey_4(57) WHEN out0_76 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_4(58) WHEN out0_76 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_4(59) WHEN out0_76 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_4(60) WHEN out0_76 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_4(61) WHEN out0_76 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_4(62) WHEN out0_76 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_4(63) WHEN out0_76 = to_unsigned(16#40#, 8) ELSE
      expandedKey_4(64) WHEN out0_76 = to_unsigned(16#41#, 8) ELSE
      expandedKey_4(65) WHEN out0_76 = to_unsigned(16#42#, 8) ELSE
      expandedKey_4(66) WHEN out0_76 = to_unsigned(16#43#, 8) ELSE
      expandedKey_4(67) WHEN out0_76 = to_unsigned(16#44#, 8) ELSE
      expandedKey_4(68) WHEN out0_76 = to_unsigned(16#45#, 8) ELSE
      expandedKey_4(69) WHEN out0_76 = to_unsigned(16#46#, 8) ELSE
      expandedKey_4(70) WHEN out0_76 = to_unsigned(16#47#, 8) ELSE
      expandedKey_4(71) WHEN out0_76 = to_unsigned(16#48#, 8) ELSE
      expandedKey_4(72) WHEN out0_76 = to_unsigned(16#49#, 8) ELSE
      expandedKey_4(73) WHEN out0_76 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_4(74) WHEN out0_76 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_4(75) WHEN out0_76 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_4(76) WHEN out0_76 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_4(77) WHEN out0_76 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_4(78) WHEN out0_76 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_4(79) WHEN out0_76 = to_unsigned(16#50#, 8) ELSE
      expandedKey_4(80) WHEN out0_76 = to_unsigned(16#51#, 8) ELSE
      expandedKey_4(81) WHEN out0_76 = to_unsigned(16#52#, 8) ELSE
      expandedKey_4(82) WHEN out0_76 = to_unsigned(16#53#, 8) ELSE
      expandedKey_4(83) WHEN out0_76 = to_unsigned(16#54#, 8) ELSE
      expandedKey_4(84) WHEN out0_76 = to_unsigned(16#55#, 8) ELSE
      expandedKey_4(85) WHEN out0_76 = to_unsigned(16#56#, 8) ELSE
      expandedKey_4(86) WHEN out0_76 = to_unsigned(16#57#, 8) ELSE
      expandedKey_4(87) WHEN out0_76 = to_unsigned(16#58#, 8) ELSE
      expandedKey_4(88) WHEN out0_76 = to_unsigned(16#59#, 8) ELSE
      expandedKey_4(89) WHEN out0_76 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_4(90) WHEN out0_76 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_4(91) WHEN out0_76 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_4(92) WHEN out0_76 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_4(93) WHEN out0_76 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_4(94) WHEN out0_76 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_4(95) WHEN out0_76 = to_unsigned(16#60#, 8) ELSE
      expandedKey_4(96) WHEN out0_76 = to_unsigned(16#61#, 8) ELSE
      expandedKey_4(97) WHEN out0_76 = to_unsigned(16#62#, 8) ELSE
      expandedKey_4(98) WHEN out0_76 = to_unsigned(16#63#, 8) ELSE
      expandedKey_4(99) WHEN out0_76 = to_unsigned(16#64#, 8) ELSE
      expandedKey_4(100) WHEN out0_76 = to_unsigned(16#65#, 8) ELSE
      expandedKey_4(101) WHEN out0_76 = to_unsigned(16#66#, 8) ELSE
      expandedKey_4(102) WHEN out0_76 = to_unsigned(16#67#, 8) ELSE
      expandedKey_4(103) WHEN out0_76 = to_unsigned(16#68#, 8) ELSE
      expandedKey_4(104) WHEN out0_76 = to_unsigned(16#69#, 8) ELSE
      expandedKey_4(105) WHEN out0_76 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_4(106) WHEN out0_76 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_4(107) WHEN out0_76 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_4(108) WHEN out0_76 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_4(109) WHEN out0_76 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_4(110) WHEN out0_76 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_4(111) WHEN out0_76 = to_unsigned(16#70#, 8) ELSE
      expandedKey_4(112) WHEN out0_76 = to_unsigned(16#71#, 8) ELSE
      expandedKey_4(113) WHEN out0_76 = to_unsigned(16#72#, 8) ELSE
      expandedKey_4(114) WHEN out0_76 = to_unsigned(16#73#, 8) ELSE
      expandedKey_4(115) WHEN out0_76 = to_unsigned(16#74#, 8) ELSE
      expandedKey_4(116) WHEN out0_76 = to_unsigned(16#75#, 8) ELSE
      expandedKey_4(117) WHEN out0_76 = to_unsigned(16#76#, 8) ELSE
      expandedKey_4(118) WHEN out0_76 = to_unsigned(16#77#, 8) ELSE
      expandedKey_4(119) WHEN out0_76 = to_unsigned(16#78#, 8) ELSE
      expandedKey_4(120) WHEN out0_76 = to_unsigned(16#79#, 8) ELSE
      expandedKey_4(121) WHEN out0_76 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_4(122) WHEN out0_76 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_4(123) WHEN out0_76 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_4(124) WHEN out0_76 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_4(125) WHEN out0_76 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_4(126) WHEN out0_76 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_4(127) WHEN out0_76 = to_unsigned(16#80#, 8) ELSE
      expandedKey_4(128) WHEN out0_76 = to_unsigned(16#81#, 8) ELSE
      expandedKey_4(129) WHEN out0_76 = to_unsigned(16#82#, 8) ELSE
      expandedKey_4(130) WHEN out0_76 = to_unsigned(16#83#, 8) ELSE
      expandedKey_4(131) WHEN out0_76 = to_unsigned(16#84#, 8) ELSE
      expandedKey_4(132) WHEN out0_76 = to_unsigned(16#85#, 8) ELSE
      expandedKey_4(133) WHEN out0_76 = to_unsigned(16#86#, 8) ELSE
      expandedKey_4(134) WHEN out0_76 = to_unsigned(16#87#, 8) ELSE
      expandedKey_4(135) WHEN out0_76 = to_unsigned(16#88#, 8) ELSE
      expandedKey_4(136) WHEN out0_76 = to_unsigned(16#89#, 8) ELSE
      expandedKey_4(137) WHEN out0_76 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_4(138) WHEN out0_76 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_4(139) WHEN out0_76 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_4(140) WHEN out0_76 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_4(141) WHEN out0_76 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_4(142) WHEN out0_76 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_4(143) WHEN out0_76 = to_unsigned(16#90#, 8) ELSE
      expandedKey_4(144) WHEN out0_76 = to_unsigned(16#91#, 8) ELSE
      expandedKey_4(145) WHEN out0_76 = to_unsigned(16#92#, 8) ELSE
      expandedKey_4(146) WHEN out0_76 = to_unsigned(16#93#, 8) ELSE
      expandedKey_4(147) WHEN out0_76 = to_unsigned(16#94#, 8) ELSE
      expandedKey_4(148) WHEN out0_76 = to_unsigned(16#95#, 8) ELSE
      expandedKey_4(149) WHEN out0_76 = to_unsigned(16#96#, 8) ELSE
      expandedKey_4(150) WHEN out0_76 = to_unsigned(16#97#, 8) ELSE
      expandedKey_4(151) WHEN out0_76 = to_unsigned(16#98#, 8) ELSE
      expandedKey_4(152) WHEN out0_76 = to_unsigned(16#99#, 8) ELSE
      expandedKey_4(153) WHEN out0_76 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_4(154) WHEN out0_76 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_4(155) WHEN out0_76 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_4(156) WHEN out0_76 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_4(157) WHEN out0_76 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_4(158) WHEN out0_76 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_4(159) WHEN out0_76 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_4(160) WHEN out0_76 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_4(161) WHEN out0_76 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_4(162) WHEN out0_76 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_4(163) WHEN out0_76 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_4(164) WHEN out0_76 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_4(165) WHEN out0_76 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_4(166) WHEN out0_76 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_4(167) WHEN out0_76 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_4(168) WHEN out0_76 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_4(169) WHEN out0_76 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_4(170) WHEN out0_76 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_4(171) WHEN out0_76 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_4(172) WHEN out0_76 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_4(173) WHEN out0_76 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_4(174) WHEN out0_76 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_4(175) WHEN out0_76 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_4(176) WHEN out0_76 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_4(177) WHEN out0_76 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_4(178) WHEN out0_76 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_4(179) WHEN out0_76 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_4(180) WHEN out0_76 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_4(181) WHEN out0_76 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_4(182) WHEN out0_76 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_4(183) WHEN out0_76 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_4(184) WHEN out0_76 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_4(185) WHEN out0_76 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_4(186) WHEN out0_76 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_4(187) WHEN out0_76 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_4(188) WHEN out0_76 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_4(189) WHEN out0_76 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_4(190) WHEN out0_76 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_4(191) WHEN out0_76 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_4(192) WHEN out0_76 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_4(193) WHEN out0_76 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_4(194) WHEN out0_76 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_4(195) WHEN out0_76 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_4(196) WHEN out0_76 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_4(197) WHEN out0_76 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_4(198) WHEN out0_76 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_4(199) WHEN out0_76 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_4(200) WHEN out0_76 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_4(201) WHEN out0_76 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_4(202) WHEN out0_76 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_4(203) WHEN out0_76 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_4(204) WHEN out0_76 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_4(205) WHEN out0_76 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_4(206) WHEN out0_76 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_4(207) WHEN out0_76 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_4(208) WHEN out0_76 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_4(209) WHEN out0_76 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_4(210) WHEN out0_76 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_4(211) WHEN out0_76 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_4(212) WHEN out0_76 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_4(213) WHEN out0_76 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_4(214) WHEN out0_76 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_4(215) WHEN out0_76 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_4(216) WHEN out0_76 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_4(217) WHEN out0_76 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_4(218) WHEN out0_76 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_4(219) WHEN out0_76 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_4(220) WHEN out0_76 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_4(221) WHEN out0_76 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_4(222) WHEN out0_76 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_4(223) WHEN out0_76 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_4(224) WHEN out0_76 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_4(225) WHEN out0_76 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_4(226) WHEN out0_76 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_4(227) WHEN out0_76 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_4(228) WHEN out0_76 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_4(229) WHEN out0_76 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_4(230) WHEN out0_76 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_4(231) WHEN out0_76 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_4(232) WHEN out0_76 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_4(233) WHEN out0_76 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_4(234) WHEN out0_76 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_4(235) WHEN out0_76 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_4(236) WHEN out0_76 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_4(237) WHEN out0_76 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_4(238) WHEN out0_76 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_4(239);

  out0_87 <= out0_86 XOR temp_key_1;

  out0_3_1 <= out0_88(3);

  
  k1_3 <= sbox(0) WHEN out0_3_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_3_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_3_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_3_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_3_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_3_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_3_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_3_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_3_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_3_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_3_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_3_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_3_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_3_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_3_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_3_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_3_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_3_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_3_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_3_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_3_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_3_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_3_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_3_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_3_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_3_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_3_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_3_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_3_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_3_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_3_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_3_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_3_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_3_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_3_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_3_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_3_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_3_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_3_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_3_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_3_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_3_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_3_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_3_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_3_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_3_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_3_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_3_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_3_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_3_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_3_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_3_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_3_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_3_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_3_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_3_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_3_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_3_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_3_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_3_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_3_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_3_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_3_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_3_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_3_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_3_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_3_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_3_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_3_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_3_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_3_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_3_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_3_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_3_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_3_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_3_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_3_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_3_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_3_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_3_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_3_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_3_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_3_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_3_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_3_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_3_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_3_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_3_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_3_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_3_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_3_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_3_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_3_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_3_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_3_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_3_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_3_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_3_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_3_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_3_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_3_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_3_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_3_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_3_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_3_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_3_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_3_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_3_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_3_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_3_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_3_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_3_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_3_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_3_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_3_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_3_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_3_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_3_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_3_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_3_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_3_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_3_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_3_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_3_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_3_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_3_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_3_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_3_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_3_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_3_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_3_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_3_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_3_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_3_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_3_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_3_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_3_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_3_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_3_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_3_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_3_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_3_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_3_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_3_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_3_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_3_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_3_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_3_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_3_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_3_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_3_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_3_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_3_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_3_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_3_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_3_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_3_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_3_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_3_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_3_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_3_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_3_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_3_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_3_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_3_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_3_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_3_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_3_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_3_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_3_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_3_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_3_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_3_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_3_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_3_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_3_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_3_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_3_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_3_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_3_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_3_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_3_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_3_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_3_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_3_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_3_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_3_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_3_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_3_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_3_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_3_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_3_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_3_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_3_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_3_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_3_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_3_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_3_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_3_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_3_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_3_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_3_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_3_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_3_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_3_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_3_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_3_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_3_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_3_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_3_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_3_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_3_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_3_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_3_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_3_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_3_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_3_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_3_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_3_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_3_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_3_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_3_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_3_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_3_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_3_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_3_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_3_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_3_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_3_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_3_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_3_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_3_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_3_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_3_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_3_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_3_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_3_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_3_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_3_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_3_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_3_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_3_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_3_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_3_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_3_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_3_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_3_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_3_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_3_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_3_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_3_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_3_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_3_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_3_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_3_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_2_1 <= out0_88(2);

  
  k1_2 <= sbox(0) WHEN out0_2_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_2_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_2_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_2_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_2_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_2_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_2_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_2_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_2_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_2_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_2_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_2_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_2_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_2_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_2_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_2_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_2_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_2_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_2_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_2_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_2_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_2_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_2_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_2_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_2_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_2_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_2_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_2_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_2_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_2_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_2_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_2_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_2_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_2_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_2_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_2_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_2_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_2_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_2_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_2_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_2_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_2_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_2_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_2_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_2_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_2_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_2_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_2_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_2_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_2_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_2_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_2_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_2_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_2_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_2_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_2_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_2_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_2_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_2_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_2_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_2_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_2_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_2_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_2_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_2_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_2_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_2_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_2_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_2_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_2_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_2_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_2_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_2_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_2_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_2_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_2_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_2_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_2_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_2_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_2_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_2_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_2_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_2_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_2_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_2_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_2_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_2_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_2_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_2_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_2_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_2_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_2_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_2_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_2_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_2_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_2_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_2_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_2_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_2_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_2_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_2_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_2_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_2_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_2_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_2_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_2_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_2_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_2_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_2_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_2_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_2_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_2_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_2_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_2_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_2_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_2_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_2_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_2_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_2_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_2_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_2_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_2_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_2_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_2_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_2_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_2_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_2_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_2_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_2_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_2_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_2_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_2_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_2_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_2_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_2_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_2_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_2_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_2_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_2_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_2_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_2_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_2_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_2_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_2_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_2_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_2_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_2_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_2_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_2_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_2_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_2_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_2_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_2_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_2_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_2_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_2_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_2_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_2_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_2_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_2_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_2_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_2_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_2_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_2_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_2_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_2_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_2_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_2_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_2_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_2_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_2_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_2_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_2_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_2_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_2_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_2_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_2_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_2_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_2_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_2_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_2_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_2_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_2_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_2_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_2_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_2_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_2_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_2_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_2_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_2_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_2_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_2_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_2_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_2_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_2_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_2_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_2_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_2_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_2_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_2_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_2_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_2_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_2_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_2_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_2_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_2_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_2_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_2_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_2_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_2_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_2_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_2_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_2_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_2_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_2_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_2_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_2_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_2_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_2_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_2_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_2_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_2_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_2_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_2_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_2_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_2_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_2_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_2_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_2_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_2_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_2_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_2_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_2_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_2_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_2_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_2_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_2_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_2_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_2_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_2_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_2_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_2_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_2_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_2_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_2_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_2_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_2_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_2_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_2_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_2_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_2_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_2_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_2_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_2_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_2_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_1_1 <= out0_88(1);

  
  k1_1 <= sbox(0) WHEN out0_1_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_1_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_1_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_1_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_1_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_1_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_1_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_1_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_1_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_1_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_1_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_1_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_1_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_1_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_1_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_1_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_1_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_1_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_1_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_1_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_1_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_1_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_1_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_1_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_1_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_1_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_1_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_1_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_1_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_1_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_1_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_1_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_1_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_1_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_1_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_1_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_1_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_1_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_1_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_1_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_1_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_1_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_1_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_1_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_1_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_1_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_1_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_1_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_1_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_1_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_1_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_1_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_1_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_1_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_1_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_1_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_1_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_1_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_1_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_1_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_1_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_1_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_1_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_1_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_1_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_1_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_1_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_1_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_1_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_1_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_1_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_1_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_1_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_1_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_1_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_1_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_1_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_1_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_1_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_1_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_1_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_1_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_1_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_1_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_1_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_1_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_1_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_1_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_1_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_1_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_1_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_1_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_1_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_1_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_1_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_1_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_1_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_1_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_1_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_1_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_1_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_1_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_1_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_1_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_1_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_1_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_1_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_1_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_1_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_1_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_1_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_1_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_1_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_1_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_1_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_1_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_1_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_1_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_1_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_1_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_1_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_1_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_1_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_1_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_1_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_1_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_1_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_1_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_1_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_1_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_1_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_1_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_1_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_1_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_1_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_1_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_1_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_1_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_1_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_1_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_1_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_1_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_1_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_1_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_1_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_1_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_1_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_1_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_1_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_1_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_1_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_1_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_1_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_1_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_1_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_1_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_1_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_1_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_1_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_1_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_1_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_1_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_1_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_1_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_1_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_1_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_1_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_1_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_1_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_1_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_1_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_1_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_1_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_1_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_1_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_1_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_1_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_1_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_1_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_1_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_1_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_1_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_1_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_1_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_1_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_1_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_1_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_1_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_1_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_1_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_1_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_1_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_1_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_1_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_1_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_1_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_1_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_1_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_1_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_1_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_1_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_1_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_1_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_1_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_1_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_1_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_1_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_1_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_1_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_1_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_1_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_1_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_1_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_1_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_1_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_1_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_1_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_1_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_1_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_1_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_1_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_1_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_1_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_1_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_1_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_1_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_1_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_1_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_1_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_1_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_1_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_1_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_1_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_1_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_1_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_1_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_1_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_1_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_1_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_1_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_1_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_1_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_1_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_1_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_1_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_1_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_1_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_1_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_1_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_1_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_1_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_1_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_1_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_1_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_1_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  rotated_key(0) <= temp_key_4(1);
  rotated_key(1) <= temp_key_4(2);
  rotated_key(2) <= temp_key_4(3);
  rotated_key(3) <= temp_key_4(0);

  out0_89(0) <= resize(rotated_key(0), 16);
  out0_89(1) <= resize(rotated_key(1), 16);
  out0_89(2) <= resize(rotated_key(2), 16);
  out0_89(3) <= resize(rotated_key(3), 16);

  out0_88(0) <= out0_89(0) + const_expression_14;
  out0_88(1) <= out0_89(1) + const_expression_14;
  out0_88(2) <= out0_89(2) + const_expression_14;
  out0_88(3) <= out0_89(3) + const_expression_14;

  out0_0 <= out0_88(0);

  
  k1_0 <= sbox(0) WHEN out0_0 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_0 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_0 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_0 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_0 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_0 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_0 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_0 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_0 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_0 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_0 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_0 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_0 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_0 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_0 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_0 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_0 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_0 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_0 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_0 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_0 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_0 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_0 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_0 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_0 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_0 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_0 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_0 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_0 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_0 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_0 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_0 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_0 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_0 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_0 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_0 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_0 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_0 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_0 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_0 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_0 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_0 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_0 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_0 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_0 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_0 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_0 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_0 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_0 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_0 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_0 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_0 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_0 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_0 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_0 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_0 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_0 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_0 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_0 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_0 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_0 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_0 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_0 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_0 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_0 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_0 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_0 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_0 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_0 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_0 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_0 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_0 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_0 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_0 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_0 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_0 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_0 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_0 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_0 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_0 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_0 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_0 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_0 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_0 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_0 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_0 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_0 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_0 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_0 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_0 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_0 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_0 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_0 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_0 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_0 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_0 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_0 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_0 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_0 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_0 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_0 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_0 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_0 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_0 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_0 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_0 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_0 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_0 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_0 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_0 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_0 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_0 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_0 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_0 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_0 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_0 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_0 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_0 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_0 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_0 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_0 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_0 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_0 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_0 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_0 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_0 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_0 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_0 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_0 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_0 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_0 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_0 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_0 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_0 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_0 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_0 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_0 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_0 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_0 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_0 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_0 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_0 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_0 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_0 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_0 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_0 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_0 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_0 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_0 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_0 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_0 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_0 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_0 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_0 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_0 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_0 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_0 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_0 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_0 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_0 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_0 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_0 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_0 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_0 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_0 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_0 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_0 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_0 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_0 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_0 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_0 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_0 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_0 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_0 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_0 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_0 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_0 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_0 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_0 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_0 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_0 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_0 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_0 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_0 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_0 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_0 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_0 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_0 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_0 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_0 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_0 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_0 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_0 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_0 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_0 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_0 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_0 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_0 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_0 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_0 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_0 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_0 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_0 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_0 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_0 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_0 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_0 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_0 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_0 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_0 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_0 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_0 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_0 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_0 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_0 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_0 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_0 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_0 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_0 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_0 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_0 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_0 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_0 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_0 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_0 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_0 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_0 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_0 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_0 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_0 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_0 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_0 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_0 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_0 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_0 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_0 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_0 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_0 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_0 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_0 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_0 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_0 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_0 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_0 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_0 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_0 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_0 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_0 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_0 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_0 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_0 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_0 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_0 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_0 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_0 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  k1(0) <= k1_0;
  k1(1) <= k1_1;
  k1(2) <= k1_2;
  k1(3) <= k1_3;

  temp_key_5(0) <= k1(0) XOR k2_1(0);
  temp_key_5(1) <= k1(1) XOR k2_1(1);
  temp_key_5(2) <= k1(2) XOR k2_1(2);
  temp_key_5(3) <= k1(3) XOR k2_1(3);

  out0_3_2 <= out0_90(3);

  
  temp_key_3_1 <= sbox(0) WHEN out0_3_2 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_3_2 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_3_2 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_3_2 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_3_2 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_3_2 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_3_2 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_3_2 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_3_2 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_3_2 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_3_2 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_3_2 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_3_2 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_3_2 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_3_2 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_3_2 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_3_2 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_3_2 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_3_2 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_3_2 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_3_2 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_3_2 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_3_2 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_3_2 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_3_2 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_3_2 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_3_2 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_3_2 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_3_2 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_3_2 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_3_2 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_3_2 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_3_2 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_3_2 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_3_2 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_3_2 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_3_2 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_3_2 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_3_2 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_3_2 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_3_2 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_3_2 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_3_2 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_3_2 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_3_2 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_3_2 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_3_2 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_3_2 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_3_2 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_3_2 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_3_2 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_3_2 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_3_2 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_3_2 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_3_2 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_3_2 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_3_2 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_3_2 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_3_2 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_3_2 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_3_2 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_3_2 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_3_2 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_3_2 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_3_2 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_3_2 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_3_2 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_3_2 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_3_2 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_3_2 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_3_2 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_3_2 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_3_2 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_3_2 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_3_2 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_3_2 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_3_2 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_3_2 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_3_2 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_3_2 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_3_2 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_3_2 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_3_2 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_3_2 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_3_2 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_3_2 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_3_2 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_3_2 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_3_2 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_3_2 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_3_2 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_3_2 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_3_2 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_3_2 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_3_2 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_3_2 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_3_2 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_3_2 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_3_2 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_3_2 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_3_2 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_3_2 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_3_2 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_3_2 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_3_2 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_3_2 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_3_2 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_3_2 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_3_2 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_3_2 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_3_2 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_3_2 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_3_2 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_3_2 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_3_2 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_3_2 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_3_2 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_3_2 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_3_2 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_3_2 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_3_2 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_3_2 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_3_2 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_3_2 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_3_2 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_3_2 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_3_2 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_3_2 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_3_2 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_3_2 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_3_2 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_3_2 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_3_2 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_3_2 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_3_2 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_3_2 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_3_2 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_3_2 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_3_2 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_3_2 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_3_2 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_3_2 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_3_2 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_3_2 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_3_2 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_3_2 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_3_2 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_3_2 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_3_2 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_3_2 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_3_2 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_3_2 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_3_2 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_3_2 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_3_2 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_3_2 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_3_2 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_3_2 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_3_2 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_3_2 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_3_2 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_3_2 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_3_2 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_3_2 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_3_2 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_3_2 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_3_2 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_3_2 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_3_2 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_3_2 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_3_2 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_3_2 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_3_2 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_3_2 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_3_2 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_3_2 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_3_2 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_3_2 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_3_2 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_3_2 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_3_2 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_3_2 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_3_2 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_3_2 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_3_2 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_3_2 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_3_2 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_3_2 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_3_2 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_3_2 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_3_2 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_3_2 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_3_2 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_3_2 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_3_2 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_3_2 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_3_2 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_3_2 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_3_2 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_3_2 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_3_2 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_3_2 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_3_2 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_3_2 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_3_2 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_3_2 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_3_2 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_3_2 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_3_2 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_3_2 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_3_2 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_3_2 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_3_2 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_3_2 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_3_2 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_3_2 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_3_2 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_3_2 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_3_2 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_3_2 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_3_2 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_3_2 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_3_2 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_3_2 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_3_2 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_3_2 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_3_2 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_3_2 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_3_2 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_3_2 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_3_2 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_3_2 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_3_2 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_3_2 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_3_2 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_3_2 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_3_2 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_3_2 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_3_2 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_3_2 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_3_2 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_3_2 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_3_2 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_3_2 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_3_2 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_3_2 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_3_2 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_3_2 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_3_2 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_3_2 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_3_2 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_3_2 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_3_2 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_3_2 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_3_2 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_2_2 <= out0_90(2);

  
  temp_key_2_1 <= sbox(0) WHEN out0_2_2 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_2_2 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_2_2 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_2_2 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_2_2 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_2_2 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_2_2 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_2_2 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_2_2 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_2_2 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_2_2 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_2_2 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_2_2 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_2_2 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_2_2 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_2_2 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_2_2 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_2_2 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_2_2 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_2_2 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_2_2 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_2_2 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_2_2 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_2_2 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_2_2 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_2_2 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_2_2 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_2_2 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_2_2 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_2_2 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_2_2 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_2_2 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_2_2 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_2_2 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_2_2 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_2_2 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_2_2 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_2_2 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_2_2 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_2_2 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_2_2 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_2_2 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_2_2 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_2_2 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_2_2 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_2_2 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_2_2 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_2_2 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_2_2 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_2_2 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_2_2 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_2_2 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_2_2 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_2_2 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_2_2 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_2_2 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_2_2 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_2_2 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_2_2 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_2_2 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_2_2 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_2_2 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_2_2 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_2_2 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_2_2 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_2_2 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_2_2 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_2_2 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_2_2 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_2_2 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_2_2 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_2_2 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_2_2 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_2_2 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_2_2 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_2_2 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_2_2 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_2_2 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_2_2 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_2_2 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_2_2 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_2_2 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_2_2 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_2_2 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_2_2 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_2_2 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_2_2 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_2_2 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_2_2 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_2_2 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_2_2 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_2_2 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_2_2 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_2_2 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_2_2 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_2_2 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_2_2 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_2_2 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_2_2 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_2_2 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_2_2 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_2_2 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_2_2 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_2_2 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_2_2 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_2_2 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_2_2 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_2_2 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_2_2 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_2_2 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_2_2 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_2_2 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_2_2 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_2_2 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_2_2 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_2_2 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_2_2 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_2_2 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_2_2 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_2_2 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_2_2 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_2_2 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_2_2 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_2_2 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_2_2 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_2_2 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_2_2 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_2_2 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_2_2 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_2_2 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_2_2 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_2_2 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_2_2 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_2_2 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_2_2 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_2_2 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_2_2 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_2_2 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_2_2 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_2_2 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_2_2 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_2_2 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_2_2 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_2_2 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_2_2 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_2_2 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_2_2 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_2_2 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_2_2 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_2_2 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_2_2 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_2_2 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_2_2 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_2_2 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_2_2 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_2_2 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_2_2 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_2_2 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_2_2 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_2_2 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_2_2 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_2_2 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_2_2 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_2_2 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_2_2 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_2_2 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_2_2 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_2_2 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_2_2 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_2_2 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_2_2 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_2_2 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_2_2 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_2_2 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_2_2 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_2_2 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_2_2 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_2_2 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_2_2 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_2_2 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_2_2 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_2_2 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_2_2 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_2_2 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_2_2 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_2_2 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_2_2 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_2_2 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_2_2 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_2_2 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_2_2 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_2_2 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_2_2 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_2_2 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_2_2 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_2_2 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_2_2 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_2_2 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_2_2 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_2_2 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_2_2 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_2_2 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_2_2 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_2_2 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_2_2 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_2_2 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_2_2 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_2_2 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_2_2 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_2_2 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_2_2 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_2_2 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_2_2 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_2_2 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_2_2 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_2_2 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_2_2 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_2_2 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_2_2 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_2_2 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_2_2 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_2_2 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_2_2 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_2_2 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_2_2 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_2_2 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_2_2 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_2_2 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_2_2 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_2_2 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_2_2 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_2_2 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_2_2 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_2_2 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_2_2 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_2_2 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_2_2 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_2_2 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_2_2 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_2_2 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_2_2 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_2_2 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_2_2 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_2_2 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_2_2 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_2_2 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_2_2 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_2_2 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_2_2 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_2_2 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_2_2 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_2_2 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_2_2 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_2_2 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_2_2 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_1_2 <= out0_90(1);

  
  temp_key_1_1 <= sbox(0) WHEN out0_1_2 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_1_2 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_1_2 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_1_2 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_1_2 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_1_2 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_1_2 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_1_2 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_1_2 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_1_2 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_1_2 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_1_2 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_1_2 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_1_2 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_1_2 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_1_2 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_1_2 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_1_2 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_1_2 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_1_2 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_1_2 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_1_2 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_1_2 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_1_2 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_1_2 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_1_2 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_1_2 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_1_2 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_1_2 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_1_2 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_1_2 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_1_2 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_1_2 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_1_2 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_1_2 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_1_2 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_1_2 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_1_2 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_1_2 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_1_2 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_1_2 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_1_2 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_1_2 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_1_2 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_1_2 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_1_2 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_1_2 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_1_2 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_1_2 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_1_2 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_1_2 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_1_2 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_1_2 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_1_2 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_1_2 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_1_2 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_1_2 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_1_2 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_1_2 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_1_2 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_1_2 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_1_2 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_1_2 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_1_2 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_1_2 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_1_2 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_1_2 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_1_2 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_1_2 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_1_2 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_1_2 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_1_2 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_1_2 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_1_2 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_1_2 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_1_2 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_1_2 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_1_2 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_1_2 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_1_2 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_1_2 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_1_2 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_1_2 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_1_2 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_1_2 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_1_2 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_1_2 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_1_2 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_1_2 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_1_2 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_1_2 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_1_2 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_1_2 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_1_2 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_1_2 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_1_2 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_1_2 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_1_2 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_1_2 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_1_2 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_1_2 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_1_2 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_1_2 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_1_2 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_1_2 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_1_2 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_1_2 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_1_2 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_1_2 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_1_2 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_1_2 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_1_2 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_1_2 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_1_2 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_1_2 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_1_2 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_1_2 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_1_2 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_1_2 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_1_2 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_1_2 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_1_2 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_1_2 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_1_2 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_1_2 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_1_2 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_1_2 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_1_2 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_1_2 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_1_2 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_1_2 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_1_2 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_1_2 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_1_2 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_1_2 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_1_2 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_1_2 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_1_2 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_1_2 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_1_2 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_1_2 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_1_2 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_1_2 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_1_2 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_1_2 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_1_2 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_1_2 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_1_2 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_1_2 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_1_2 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_1_2 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_1_2 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_1_2 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_1_2 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_1_2 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_1_2 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_1_2 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_1_2 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_1_2 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_1_2 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_1_2 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_1_2 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_1_2 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_1_2 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_1_2 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_1_2 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_1_2 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_1_2 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_1_2 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_1_2 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_1_2 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_1_2 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_1_2 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_1_2 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_1_2 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_1_2 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_1_2 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_1_2 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_1_2 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_1_2 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_1_2 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_1_2 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_1_2 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_1_2 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_1_2 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_1_2 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_1_2 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_1_2 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_1_2 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_1_2 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_1_2 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_1_2 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_1_2 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_1_2 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_1_2 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_1_2 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_1_2 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_1_2 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_1_2 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_1_2 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_1_2 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_1_2 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_1_2 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_1_2 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_1_2 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_1_2 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_1_2 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_1_2 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_1_2 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_1_2 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_1_2 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_1_2 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_1_2 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_1_2 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_1_2 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_1_2 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_1_2 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_1_2 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_1_2 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_1_2 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_1_2 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_1_2 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_1_2 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_1_2 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_1_2 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_1_2 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_1_2 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_1_2 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_1_2 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_1_2 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_1_2 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_1_2 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_1_2 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_1_2 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_1_2 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_1_2 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_1_2 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_1_2 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_1_2 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_1_2 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_1_2 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_1_2 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_1_2 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_1_2 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_1_2 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_1_2 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_1_2 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_1_2 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_1_2 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_1_2 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_1_2 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_1_2 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_1_2 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_1_2 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_1_2 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_91(0) <= resize(temp_key_4(0), 16);
  out0_91(1) <= resize(temp_key_4(1), 16);
  out0_91(2) <= resize(temp_key_4(2), 16);
  out0_91(3) <= resize(temp_key_4(3), 16);

  out0_90(0) <= out0_91(0) + const_expression_13;
  out0_90(1) <= out0_91(1) + const_expression_13;
  out0_90(2) <= out0_91(2) + const_expression_13;
  out0_90(3) <= out0_91(3) + const_expression_13;

  out0_0_1 <= out0_90(0);

  
  temp_key_0 <= sbox(0) WHEN out0_0_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_0_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_0_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_0_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_0_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_0_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_0_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_0_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_0_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_0_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_0_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_0_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_0_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_0_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_0_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_0_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_0_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_0_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_0_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_0_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_0_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_0_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_0_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_0_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_0_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_0_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_0_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_0_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_0_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_0_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_0_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_0_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_0_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_0_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_0_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_0_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_0_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_0_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_0_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_0_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_0_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_0_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_0_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_0_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_0_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_0_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_0_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_0_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_0_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_0_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_0_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_0_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_0_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_0_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_0_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_0_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_0_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_0_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_0_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_0_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_0_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_0_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_0_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_0_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_0_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_0_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_0_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_0_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_0_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_0_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_0_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_0_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_0_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_0_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_0_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_0_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_0_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_0_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_0_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_0_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_0_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_0_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_0_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_0_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_0_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_0_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_0_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_0_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_0_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_0_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_0_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_0_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_0_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_0_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_0_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_0_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_0_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_0_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_0_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_0_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_0_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_0_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_0_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_0_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_0_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_0_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_0_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_0_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_0_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_0_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_0_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_0_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_0_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_0_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_0_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_0_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_0_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_0_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_0_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_0_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_0_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_0_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_0_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_0_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_0_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_0_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_0_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_0_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_0_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_0_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_0_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_0_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_0_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_0_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_0_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_0_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_0_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_0_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_0_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_0_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_0_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_0_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_0_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_0_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_0_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_0_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_0_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_0_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_0_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_0_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_0_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_0_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_0_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_0_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_0_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_0_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_0_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_0_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_0_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_0_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_0_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_0_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_0_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_0_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_0_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_0_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_0_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_0_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_0_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_0_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_0_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_0_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_0_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_0_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_0_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_0_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_0_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_0_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_0_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_0_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_0_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_0_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_0_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_0_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_0_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_0_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_0_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_0_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_0_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_0_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_0_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_0_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_0_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_0_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_0_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_0_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_0_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_0_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_0_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_0_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_0_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_0_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_0_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_0_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_0_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_0_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_0_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_0_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_0_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_0_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_0_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_0_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_0_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_0_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_0_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_0_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_0_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_0_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_0_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_0_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_0_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_0_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_0_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_0_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_0_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_0_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_0_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_0_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_0_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_0_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_0_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_0_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_0_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_0_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_0_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_0_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_0_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_0_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_0_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_0_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_0_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_0_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_0_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_0_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_0_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_0_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_0_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_0_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_0_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_0_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_0_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_0_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_0_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_0_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_0_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  temp_key_6(0) <= temp_key_0;
  temp_key_6(1) <= temp_key_1_1;
  temp_key_6(2) <= temp_key_2_1;
  temp_key_6(3) <= temp_key_3_1;

  
  out0_92 <= expandedKey(0) WHEN out0_54 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_54 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_54 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_54 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_54 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_54 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_54 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_54 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_54 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_54 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_54 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_54 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_54 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_54 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_54 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_54 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_54 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_54 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_54 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_54 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_54 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_54 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_54 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_54 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_54 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_54 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_54 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_54 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_54 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_54 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_54 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_54 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_54 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_54 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_54 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_54 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_54 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_54 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_54 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_54 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_54 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_54 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_54 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_54 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_54 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_54 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_54 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_54 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_54 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_54 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_54 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_54 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_54 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_54 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_54 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_54 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_54 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_54 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_54 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_54 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_54 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_54 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_54 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_54 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_54 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_54 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_54 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_54 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_54 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_54 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_54 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_54 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_54 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_54 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_54 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_54 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_54 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_54 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_54 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_54 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_54 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_54 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_54 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_54 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_54 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_54 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_54 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_54 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_54 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_54 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_54 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_54 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_54 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_54 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_54 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_54 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_54 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_54 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_54 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_54 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_54 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_54 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_54 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_54 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_54 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_54 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_54 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_54 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_54 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_54 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_54 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_54 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_54 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_54 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_54 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_54 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_54 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_54 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_54 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_54 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_54 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_54 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_54 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_54 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_54 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_54 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_54 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_54 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_54 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_54 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_54 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_54 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_54 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_54 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_54 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_54 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_54 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_54 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_54 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_54 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_54 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_54 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_54 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_54 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_54 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_54 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_54 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_54 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_54 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_54 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_54 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_54 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_54 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_54 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_54 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_54 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_54 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_54 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_54 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_54 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_54 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_54 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_54 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_54 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_54 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_54 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_54 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_54 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_54 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_54 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_54 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_54 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_54 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_54 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_54 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_54 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_54 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_54 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_54 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_54 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_54 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_54 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_54 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_54 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_54 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_54 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_54 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_54 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_54 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_54 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_54 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_54 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_54 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_54 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_54 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_54 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_54 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_54 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_54 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_54 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_54 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_54 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_54 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_54 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_54 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_54 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_54 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_54 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_54 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_54 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_54 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_54 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_54 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_54 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_54 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_54 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_54 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_54 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_54 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_54 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_54 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_54 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_54 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_54 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_54 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_54 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_54 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_54 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_54 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_54 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_54 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_54 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_54 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_54 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_54 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_54 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_54 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_54 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_54 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  
  out0_93 <= expandedKey(0) WHEN out0_53 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_53 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_53 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_53 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_53 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_53 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_53 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_53 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_53 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_53 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_53 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_53 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_53 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_53 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_53 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_53 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_53 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_53 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_53 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_53 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_53 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_53 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_53 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_53 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_53 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_53 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_53 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_53 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_53 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_53 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_53 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_53 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_53 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_53 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_53 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_53 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_53 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_53 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_53 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_53 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_53 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_53 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_53 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_53 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_53 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_53 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_53 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_53 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_53 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_53 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_53 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_53 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_53 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_53 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_53 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_53 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_53 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_53 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_53 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_53 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_53 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_53 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_53 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_53 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_53 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_53 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_53 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_53 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_53 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_53 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_53 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_53 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_53 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_53 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_53 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_53 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_53 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_53 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_53 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_53 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_53 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_53 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_53 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_53 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_53 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_53 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_53 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_53 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_53 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_53 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_53 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_53 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_53 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_53 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_53 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_53 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_53 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_53 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_53 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_53 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_53 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_53 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_53 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_53 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_53 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_53 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_53 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_53 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_53 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_53 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_53 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_53 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_53 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_53 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_53 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_53 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_53 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_53 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_53 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_53 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_53 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_53 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_53 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_53 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_53 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_53 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_53 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_53 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_53 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_53 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_53 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_53 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_53 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_53 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_53 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_53 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_53 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_53 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_53 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_53 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_53 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_53 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_53 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_53 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_53 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_53 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_53 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_53 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_53 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_53 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_53 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_53 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_53 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_53 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_53 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_53 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_53 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_53 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_53 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_53 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_53 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_53 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_53 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_53 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_53 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_53 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_53 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_53 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_53 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_53 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_53 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_53 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_53 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_53 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_53 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_53 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_53 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_53 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_53 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_53 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_53 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_53 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_53 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_53 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_53 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_53 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_53 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_53 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_53 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_53 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_53 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_53 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_53 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_53 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_53 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_53 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_53 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_53 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_53 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_53 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_53 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_53 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_53 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_53 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_53 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_53 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_53 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_53 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_53 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_53 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_53 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_53 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_53 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_53 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_53 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_53 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_53 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_53 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_53 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_53 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_53 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_53 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_53 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_53 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_53 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_53 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_53 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_53 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_53 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_53 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_53 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_53 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_53 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_53 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_53 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_53 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_53 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_53 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_53 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  
  out0_94 <= expandedKey(0) WHEN out0_52 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_52 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_52 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_52 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_52 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_52 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_52 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_52 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_52 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_52 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_52 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_52 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_52 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_52 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_52 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_52 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_52 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_52 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_52 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_52 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_52 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_52 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_52 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_52 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_52 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_52 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_52 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_52 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_52 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_52 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_52 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_52 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_52 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_52 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_52 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_52 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_52 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_52 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_52 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_52 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_52 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_52 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_52 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_52 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_52 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_52 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_52 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_52 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_52 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_52 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_52 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_52 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_52 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_52 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_52 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_52 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_52 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_52 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_52 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_52 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_52 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_52 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_52 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_52 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_52 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_52 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_52 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_52 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_52 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_52 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_52 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_52 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_52 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_52 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_52 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_52 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_52 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_52 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_52 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_52 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_52 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_52 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_52 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_52 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_52 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_52 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_52 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_52 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_52 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_52 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_52 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_52 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_52 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_52 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_52 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_52 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_52 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_52 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_52 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_52 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_52 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_52 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_52 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_52 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_52 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_52 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_52 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_52 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_52 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_52 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_52 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_52 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_52 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_52 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_52 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_52 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_52 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_52 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_52 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_52 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_52 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_52 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_52 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_52 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_52 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_52 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_52 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_52 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_52 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_52 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_52 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_52 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_52 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_52 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_52 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_52 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_52 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_52 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_52 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_52 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_52 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_52 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_52 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_52 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_52 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_52 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_52 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_52 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_52 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_52 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_52 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_52 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_52 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_52 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_52 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_52 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_52 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_52 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_52 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_52 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_52 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_52 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_52 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_52 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_52 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_52 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_52 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_52 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_52 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_52 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_52 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_52 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_52 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_52 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_52 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_52 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_52 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_52 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_52 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_52 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_52 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_52 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_52 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_52 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_52 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_52 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_52 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_52 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_52 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_52 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_52 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_52 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_52 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_52 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_52 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_52 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_52 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_52 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_52 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_52 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_52 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_52 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_52 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_52 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_52 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_52 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_52 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_52 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_52 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_52 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_52 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_52 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_52 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_52 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_52 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_52 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_52 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_52 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_52 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_52 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_52 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_52 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_52 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_52 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_52 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_52 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_52 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_52 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_52 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_52 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_52 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_52 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_52 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_52 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_52 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_52 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_52 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_52 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_52 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  
  out0_95 <= expandedKey(0) WHEN out0_51 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_51 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_51 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_51 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_51 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_51 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_51 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_51 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_51 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_51 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_51 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_51 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_51 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_51 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_51 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_51 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_51 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_51 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_51 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_51 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_51 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_51 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_51 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_51 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_51 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_51 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_51 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_51 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_51 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_51 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_51 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_51 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_51 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_51 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_51 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_51 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_51 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_51 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_51 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_51 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_51 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_51 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_51 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_51 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_51 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_51 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_51 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_51 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_51 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_51 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_51 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_51 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_51 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_51 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_51 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_51 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_51 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_51 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_51 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_51 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_51 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_51 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_51 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_51 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_51 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_51 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_51 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_51 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_51 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_51 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_51 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_51 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_51 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_51 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_51 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_51 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_51 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_51 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_51 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_51 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_51 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_51 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_51 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_51 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_51 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_51 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_51 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_51 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_51 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_51 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_51 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_51 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_51 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_51 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_51 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_51 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_51 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_51 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_51 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_51 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_51 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_51 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_51 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_51 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_51 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_51 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_51 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_51 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_51 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_51 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_51 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_51 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_51 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_51 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_51 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_51 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_51 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_51 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_51 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_51 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_51 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_51 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_51 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_51 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_51 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_51 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_51 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_51 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_51 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_51 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_51 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_51 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_51 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_51 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_51 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_51 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_51 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_51 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_51 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_51 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_51 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_51 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_51 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_51 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_51 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_51 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_51 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_51 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_51 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_51 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_51 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_51 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_51 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_51 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_51 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_51 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_51 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_51 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_51 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_51 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_51 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_51 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_51 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_51 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_51 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_51 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_51 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_51 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_51 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_51 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_51 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_51 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_51 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_51 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_51 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_51 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_51 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_51 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_51 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_51 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_51 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_51 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_51 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_51 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_51 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_51 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_51 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_51 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_51 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_51 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_51 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_51 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_51 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_51 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_51 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_51 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_51 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_51 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_51 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_51 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_51 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_51 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_51 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_51 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_51 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_51 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_51 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_51 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_51 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_51 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_51 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_51 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_51 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_51 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_51 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_51 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_51 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_51 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_51 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_51 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_51 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_51 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_51 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_51 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_51 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_51 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_51 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_51 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_51 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_51 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_51 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_51 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_51 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_51 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_51 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_51 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_51 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_51 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_51 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  
  out0_96(0) <= temp_key_7(0) WHEN out0_10 = '0' ELSE
      temp_key_7(0);
  
  out0_96(1) <= temp_key_7(1) WHEN out0_10 = '0' ELSE
      temp_key_7(1);
  
  out0_96(2) <= temp_key_7(2) WHEN out0_10 = '0' ELSE
      temp_key_7(2);
  
  out0_96(3) <= temp_key_7(3) WHEN out0_10 = '0' ELSE
      temp_key_7(3);

  
  out0_97(0) <= out0_96(0) WHEN out0_12 = '0' ELSE
      temp_key_7(0);
  
  out0_97(1) <= out0_96(1) WHEN out0_12 = '0' ELSE
      temp_key_7(1);
  
  out0_97(2) <= out0_96(2) WHEN out0_12 = '0' ELSE
      temp_key_7(2);
  
  out0_97(3) <= out0_96(3) WHEN out0_12 = '0' ELSE
      temp_key_7(3);

  
  out0_98(0) <= out0_97(0) WHEN out0_14 = '0' ELSE
      temp_key_7(0);
  
  out0_98(1) <= out0_97(1) WHEN out0_14 = '0' ELSE
      temp_key_7(1);
  
  out0_98(2) <= out0_97(2) WHEN out0_14 = '0' ELSE
      temp_key_7(2);
  
  out0_98(3) <= out0_97(3) WHEN out0_14 = '0' ELSE
      temp_key_7(3);

  
  out0_99(0) <= out0_98(0) WHEN out0_16 = '0' ELSE
      temp_key_7(0);
  
  out0_99(1) <= out0_98(1) WHEN out0_16 = '0' ELSE
      temp_key_7(1);
  
  out0_99(2) <= out0_98(2) WHEN out0_16 = '0' ELSE
      temp_key_7(2);
  
  out0_99(3) <= out0_98(3) WHEN out0_16 = '0' ELSE
      temp_key_7(3);

  
  out0_100(0) <= out0_99(0) WHEN out0_18 = '0' ELSE
      temp_key_7(0);
  
  out0_100(1) <= out0_99(1) WHEN out0_18 = '0' ELSE
      temp_key_7(1);
  
  out0_100(2) <= out0_99(2) WHEN out0_18 = '0' ELSE
      temp_key_7(2);
  
  out0_100(3) <= out0_99(3) WHEN out0_18 = '0' ELSE
      temp_key_7(3);

  
  out0_101(0) <= out0_100(0) WHEN out0_20 = '0' ELSE
      temp_key_7(0);
  
  out0_101(1) <= out0_100(1) WHEN out0_20 = '0' ELSE
      temp_key_7(1);
  
  out0_101(2) <= out0_100(2) WHEN out0_20 = '0' ELSE
      temp_key_7(2);
  
  out0_101(3) <= out0_100(3) WHEN out0_20 = '0' ELSE
      temp_key_7(3);

  
  out0_102(0) <= out0_101(0) WHEN out0_22 = '0' ELSE
      temp_key(0);
  
  out0_102(1) <= out0_101(1) WHEN out0_22 = '0' ELSE
      temp_key(1);
  
  out0_102(2) <= out0_101(2) WHEN out0_22 = '0' ELSE
      temp_key(2);
  
  out0_102(3) <= out0_101(3) WHEN out0_22 = '0' ELSE
      temp_key(3);

  
  temp_key_8(0) <= out0_102(0) WHEN out0_24 = '0' ELSE
      temp_key_7(0);
  
  temp_key_8(1) <= out0_102(1) WHEN out0_24 = '0' ELSE
      temp_key_7(1);
  
  temp_key_8(2) <= out0_102(2) WHEN out0_24 = '0' ELSE
      temp_key_7(2);
  
  temp_key_8(3) <= out0_102(3) WHEN out0_24 = '0' ELSE
      temp_key_7(3);

  intdelay9_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        temp_key_7(0) <= to_unsigned(16#00#, 8);
        temp_key_7(1) <= to_unsigned(16#00#, 8);
        temp_key_7(2) <= to_unsigned(16#00#, 8);
        temp_key_7(3) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        temp_key_7(0) <= temp_key_8(0);
        temp_key_7(1) <= temp_key_8(1);
        temp_key_7(2) <= temp_key_8(2);
        temp_key_7(3) <= temp_key_8(3);
      END IF;
    END IF;
  END PROCESS intdelay9_process;


  temp_key_9(0) <= out0_95;
  temp_key_9(1) <= temp_key_7(1);
  temp_key_9(2) <= temp_key_7(2);
  temp_key_9(3) <= temp_key_7(3);

  temp_key_10(0) <= temp_key_9(0);
  temp_key_10(1) <= out0_94;
  temp_key_10(2) <= temp_key_9(2);
  temp_key_10(3) <= temp_key_9(3);

  temp_key_11(0) <= temp_key_10(0);
  temp_key_11(1) <= temp_key_10(1);
  temp_key_11(2) <= out0_93;
  temp_key_11(3) <= temp_key_10(3);

  temp_key_4(0) <= temp_key_11(0);
  temp_key_4(1) <= temp_key_11(1);
  temp_key_4(2) <= temp_key_11(2);
  temp_key_4(3) <= out0_92;

  
  out0_103(0) <= temp_key_4(0) WHEN out0_5 = '0' ELSE
      temp_key_6(0);
  
  out0_103(1) <= temp_key_4(1) WHEN out0_5 = '0' ELSE
      temp_key_6(1);
  
  out0_103(2) <= temp_key_4(2) WHEN out0_5 = '0' ELSE
      temp_key_6(2);
  
  out0_103(3) <= temp_key_4(3) WHEN out0_5 = '0' ELSE
      temp_key_6(3);

  
  temp_key(0) <= out0_103(0) WHEN out0_9 = '0' ELSE
      temp_key_5(0);
  
  temp_key(1) <= out0_103(1) WHEN out0_9 = '0' ELSE
      temp_key_5(1);
  
  temp_key(2) <= out0_103(2) WHEN out0_9 = '0' ELSE
      temp_key_5(2);
  
  temp_key(3) <= out0_103(3) WHEN out0_9 = '0' ELSE
      temp_key_5(3);

  temp_key_0_1 <= temp_key(0);

  
  out0_104 <= expandedKey(0) WHEN out0_50 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_50 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_50 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_50 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_50 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_50 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_50 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_50 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_50 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_50 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_50 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_50 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_50 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_50 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_50 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_50 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_50 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_50 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_50 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_50 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_50 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_50 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_50 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_50 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_50 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_50 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_50 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_50 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_50 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_50 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_50 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_50 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_50 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_50 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_50 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_50 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_50 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_50 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_50 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_50 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_50 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_50 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_50 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_50 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_50 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_50 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_50 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_50 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_50 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_50 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_50 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_50 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_50 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_50 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_50 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_50 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_50 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_50 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_50 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_50 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_50 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_50 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_50 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_50 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_50 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_50 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_50 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_50 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_50 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_50 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_50 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_50 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_50 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_50 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_50 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_50 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_50 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_50 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_50 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_50 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_50 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_50 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_50 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_50 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_50 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_50 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_50 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_50 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_50 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_50 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_50 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_50 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_50 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_50 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_50 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_50 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_50 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_50 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_50 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_50 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_50 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_50 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_50 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_50 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_50 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_50 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_50 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_50 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_50 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_50 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_50 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_50 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_50 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_50 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_50 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_50 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_50 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_50 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_50 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_50 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_50 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_50 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_50 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_50 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_50 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_50 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_50 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_50 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_50 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_50 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_50 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_50 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_50 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_50 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_50 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_50 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_50 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_50 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_50 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_50 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_50 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_50 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_50 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_50 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_50 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_50 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_50 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_50 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_50 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_50 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_50 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_50 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_50 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_50 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_50 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_50 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_50 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_50 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_50 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_50 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_50 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_50 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_50 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_50 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_50 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_50 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_50 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_50 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_50 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_50 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_50 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_50 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_50 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_50 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_50 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_50 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_50 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_50 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_50 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_50 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_50 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_50 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_50 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_50 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_50 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_50 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_50 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_50 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_50 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_50 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_50 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_50 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_50 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_50 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_50 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_50 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_50 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_50 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_50 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_50 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_50 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_50 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_50 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_50 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_50 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_50 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_50 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_50 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_50 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_50 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_50 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_50 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_50 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_50 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_50 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_50 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_50 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_50 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_50 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_50 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_50 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_50 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_50 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_50 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_50 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_50 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_50 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_50 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_50 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_50 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_50 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_50 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_50 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_50 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_50 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_50 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_50 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_50 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_50 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  out0_105 <= out0_104 XOR temp_key_0_1;

  
  expandedKey_4(0) <= out0_105 WHEN out0_75 = to_unsigned(16#01#, 8) ELSE
      expandedKey(0);
  
  expandedKey_4(1) <= out0_105 WHEN out0_75 = to_unsigned(16#02#, 8) ELSE
      expandedKey(1);
  
  expandedKey_4(2) <= out0_105 WHEN out0_75 = to_unsigned(16#03#, 8) ELSE
      expandedKey(2);
  
  expandedKey_4(3) <= out0_105 WHEN out0_75 = to_unsigned(16#04#, 8) ELSE
      expandedKey(3);
  
  expandedKey_4(4) <= out0_105 WHEN out0_75 = to_unsigned(16#05#, 8) ELSE
      expandedKey(4);
  
  expandedKey_4(5) <= out0_105 WHEN out0_75 = to_unsigned(16#06#, 8) ELSE
      expandedKey(5);
  
  expandedKey_4(6) <= out0_105 WHEN out0_75 = to_unsigned(16#07#, 8) ELSE
      expandedKey(6);
  
  expandedKey_4(7) <= out0_105 WHEN out0_75 = to_unsigned(16#08#, 8) ELSE
      expandedKey(7);
  
  expandedKey_4(8) <= out0_105 WHEN out0_75 = to_unsigned(16#09#, 8) ELSE
      expandedKey(8);
  
  expandedKey_4(9) <= out0_105 WHEN out0_75 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(9);
  
  expandedKey_4(10) <= out0_105 WHEN out0_75 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(10);
  
  expandedKey_4(11) <= out0_105 WHEN out0_75 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(11);
  
  expandedKey_4(12) <= out0_105 WHEN out0_75 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(12);
  
  expandedKey_4(13) <= out0_105 WHEN out0_75 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(13);
  
  expandedKey_4(14) <= out0_105 WHEN out0_75 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(14);
  
  expandedKey_4(15) <= out0_105 WHEN out0_75 = to_unsigned(16#10#, 8) ELSE
      expandedKey(15);
  
  expandedKey_4(16) <= out0_105 WHEN out0_75 = to_unsigned(16#11#, 8) ELSE
      expandedKey(16);
  
  expandedKey_4(17) <= out0_105 WHEN out0_75 = to_unsigned(16#12#, 8) ELSE
      expandedKey(17);
  
  expandedKey_4(18) <= out0_105 WHEN out0_75 = to_unsigned(16#13#, 8) ELSE
      expandedKey(18);
  
  expandedKey_4(19) <= out0_105 WHEN out0_75 = to_unsigned(16#14#, 8) ELSE
      expandedKey(19);
  
  expandedKey_4(20) <= out0_105 WHEN out0_75 = to_unsigned(16#15#, 8) ELSE
      expandedKey(20);
  
  expandedKey_4(21) <= out0_105 WHEN out0_75 = to_unsigned(16#16#, 8) ELSE
      expandedKey(21);
  
  expandedKey_4(22) <= out0_105 WHEN out0_75 = to_unsigned(16#17#, 8) ELSE
      expandedKey(22);
  
  expandedKey_4(23) <= out0_105 WHEN out0_75 = to_unsigned(16#18#, 8) ELSE
      expandedKey(23);
  
  expandedKey_4(24) <= out0_105 WHEN out0_75 = to_unsigned(16#19#, 8) ELSE
      expandedKey(24);
  
  expandedKey_4(25) <= out0_105 WHEN out0_75 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(25);
  
  expandedKey_4(26) <= out0_105 WHEN out0_75 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(26);
  
  expandedKey_4(27) <= out0_105 WHEN out0_75 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(27);
  
  expandedKey_4(28) <= out0_105 WHEN out0_75 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(28);
  
  expandedKey_4(29) <= out0_105 WHEN out0_75 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(29);
  
  expandedKey_4(30) <= out0_105 WHEN out0_75 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(30);
  
  expandedKey_4(31) <= out0_105 WHEN out0_75 = to_unsigned(16#20#, 8) ELSE
      expandedKey(31);
  
  expandedKey_4(32) <= out0_105 WHEN out0_75 = to_unsigned(16#21#, 8) ELSE
      expandedKey(32);
  
  expandedKey_4(33) <= out0_105 WHEN out0_75 = to_unsigned(16#22#, 8) ELSE
      expandedKey(33);
  
  expandedKey_4(34) <= out0_105 WHEN out0_75 = to_unsigned(16#23#, 8) ELSE
      expandedKey(34);
  
  expandedKey_4(35) <= out0_105 WHEN out0_75 = to_unsigned(16#24#, 8) ELSE
      expandedKey(35);
  
  expandedKey_4(36) <= out0_105 WHEN out0_75 = to_unsigned(16#25#, 8) ELSE
      expandedKey(36);
  
  expandedKey_4(37) <= out0_105 WHEN out0_75 = to_unsigned(16#26#, 8) ELSE
      expandedKey(37);
  
  expandedKey_4(38) <= out0_105 WHEN out0_75 = to_unsigned(16#27#, 8) ELSE
      expandedKey(38);
  
  expandedKey_4(39) <= out0_105 WHEN out0_75 = to_unsigned(16#28#, 8) ELSE
      expandedKey(39);
  
  expandedKey_4(40) <= out0_105 WHEN out0_75 = to_unsigned(16#29#, 8) ELSE
      expandedKey(40);
  
  expandedKey_4(41) <= out0_105 WHEN out0_75 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(41);
  
  expandedKey_4(42) <= out0_105 WHEN out0_75 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(42);
  
  expandedKey_4(43) <= out0_105 WHEN out0_75 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(43);
  
  expandedKey_4(44) <= out0_105 WHEN out0_75 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(44);
  
  expandedKey_4(45) <= out0_105 WHEN out0_75 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(45);
  
  expandedKey_4(46) <= out0_105 WHEN out0_75 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(46);
  
  expandedKey_4(47) <= out0_105 WHEN out0_75 = to_unsigned(16#30#, 8) ELSE
      expandedKey(47);
  
  expandedKey_4(48) <= out0_105 WHEN out0_75 = to_unsigned(16#31#, 8) ELSE
      expandedKey(48);
  
  expandedKey_4(49) <= out0_105 WHEN out0_75 = to_unsigned(16#32#, 8) ELSE
      expandedKey(49);
  
  expandedKey_4(50) <= out0_105 WHEN out0_75 = to_unsigned(16#33#, 8) ELSE
      expandedKey(50);
  
  expandedKey_4(51) <= out0_105 WHEN out0_75 = to_unsigned(16#34#, 8) ELSE
      expandedKey(51);
  
  expandedKey_4(52) <= out0_105 WHEN out0_75 = to_unsigned(16#35#, 8) ELSE
      expandedKey(52);
  
  expandedKey_4(53) <= out0_105 WHEN out0_75 = to_unsigned(16#36#, 8) ELSE
      expandedKey(53);
  
  expandedKey_4(54) <= out0_105 WHEN out0_75 = to_unsigned(16#37#, 8) ELSE
      expandedKey(54);
  
  expandedKey_4(55) <= out0_105 WHEN out0_75 = to_unsigned(16#38#, 8) ELSE
      expandedKey(55);
  
  expandedKey_4(56) <= out0_105 WHEN out0_75 = to_unsigned(16#39#, 8) ELSE
      expandedKey(56);
  
  expandedKey_4(57) <= out0_105 WHEN out0_75 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(57);
  
  expandedKey_4(58) <= out0_105 WHEN out0_75 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(58);
  
  expandedKey_4(59) <= out0_105 WHEN out0_75 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(59);
  
  expandedKey_4(60) <= out0_105 WHEN out0_75 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(60);
  
  expandedKey_4(61) <= out0_105 WHEN out0_75 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(61);
  
  expandedKey_4(62) <= out0_105 WHEN out0_75 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(62);
  
  expandedKey_4(63) <= out0_105 WHEN out0_75 = to_unsigned(16#40#, 8) ELSE
      expandedKey(63);
  
  expandedKey_4(64) <= out0_105 WHEN out0_75 = to_unsigned(16#41#, 8) ELSE
      expandedKey(64);
  
  expandedKey_4(65) <= out0_105 WHEN out0_75 = to_unsigned(16#42#, 8) ELSE
      expandedKey(65);
  
  expandedKey_4(66) <= out0_105 WHEN out0_75 = to_unsigned(16#43#, 8) ELSE
      expandedKey(66);
  
  expandedKey_4(67) <= out0_105 WHEN out0_75 = to_unsigned(16#44#, 8) ELSE
      expandedKey(67);
  
  expandedKey_4(68) <= out0_105 WHEN out0_75 = to_unsigned(16#45#, 8) ELSE
      expandedKey(68);
  
  expandedKey_4(69) <= out0_105 WHEN out0_75 = to_unsigned(16#46#, 8) ELSE
      expandedKey(69);
  
  expandedKey_4(70) <= out0_105 WHEN out0_75 = to_unsigned(16#47#, 8) ELSE
      expandedKey(70);
  
  expandedKey_4(71) <= out0_105 WHEN out0_75 = to_unsigned(16#48#, 8) ELSE
      expandedKey(71);
  
  expandedKey_4(72) <= out0_105 WHEN out0_75 = to_unsigned(16#49#, 8) ELSE
      expandedKey(72);
  
  expandedKey_4(73) <= out0_105 WHEN out0_75 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(73);
  
  expandedKey_4(74) <= out0_105 WHEN out0_75 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(74);
  
  expandedKey_4(75) <= out0_105 WHEN out0_75 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(75);
  
  expandedKey_4(76) <= out0_105 WHEN out0_75 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(76);
  
  expandedKey_4(77) <= out0_105 WHEN out0_75 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(77);
  
  expandedKey_4(78) <= out0_105 WHEN out0_75 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(78);
  
  expandedKey_4(79) <= out0_105 WHEN out0_75 = to_unsigned(16#50#, 8) ELSE
      expandedKey(79);
  
  expandedKey_4(80) <= out0_105 WHEN out0_75 = to_unsigned(16#51#, 8) ELSE
      expandedKey(80);
  
  expandedKey_4(81) <= out0_105 WHEN out0_75 = to_unsigned(16#52#, 8) ELSE
      expandedKey(81);
  
  expandedKey_4(82) <= out0_105 WHEN out0_75 = to_unsigned(16#53#, 8) ELSE
      expandedKey(82);
  
  expandedKey_4(83) <= out0_105 WHEN out0_75 = to_unsigned(16#54#, 8) ELSE
      expandedKey(83);
  
  expandedKey_4(84) <= out0_105 WHEN out0_75 = to_unsigned(16#55#, 8) ELSE
      expandedKey(84);
  
  expandedKey_4(85) <= out0_105 WHEN out0_75 = to_unsigned(16#56#, 8) ELSE
      expandedKey(85);
  
  expandedKey_4(86) <= out0_105 WHEN out0_75 = to_unsigned(16#57#, 8) ELSE
      expandedKey(86);
  
  expandedKey_4(87) <= out0_105 WHEN out0_75 = to_unsigned(16#58#, 8) ELSE
      expandedKey(87);
  
  expandedKey_4(88) <= out0_105 WHEN out0_75 = to_unsigned(16#59#, 8) ELSE
      expandedKey(88);
  
  expandedKey_4(89) <= out0_105 WHEN out0_75 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(89);
  
  expandedKey_4(90) <= out0_105 WHEN out0_75 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(90);
  
  expandedKey_4(91) <= out0_105 WHEN out0_75 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(91);
  
  expandedKey_4(92) <= out0_105 WHEN out0_75 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(92);
  
  expandedKey_4(93) <= out0_105 WHEN out0_75 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(93);
  
  expandedKey_4(94) <= out0_105 WHEN out0_75 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(94);
  
  expandedKey_4(95) <= out0_105 WHEN out0_75 = to_unsigned(16#60#, 8) ELSE
      expandedKey(95);
  
  expandedKey_4(96) <= out0_105 WHEN out0_75 = to_unsigned(16#61#, 8) ELSE
      expandedKey(96);
  
  expandedKey_4(97) <= out0_105 WHEN out0_75 = to_unsigned(16#62#, 8) ELSE
      expandedKey(97);
  
  expandedKey_4(98) <= out0_105 WHEN out0_75 = to_unsigned(16#63#, 8) ELSE
      expandedKey(98);
  
  expandedKey_4(99) <= out0_105 WHEN out0_75 = to_unsigned(16#64#, 8) ELSE
      expandedKey(99);
  
  expandedKey_4(100) <= out0_105 WHEN out0_75 = to_unsigned(16#65#, 8) ELSE
      expandedKey(100);
  
  expandedKey_4(101) <= out0_105 WHEN out0_75 = to_unsigned(16#66#, 8) ELSE
      expandedKey(101);
  
  expandedKey_4(102) <= out0_105 WHEN out0_75 = to_unsigned(16#67#, 8) ELSE
      expandedKey(102);
  
  expandedKey_4(103) <= out0_105 WHEN out0_75 = to_unsigned(16#68#, 8) ELSE
      expandedKey(103);
  
  expandedKey_4(104) <= out0_105 WHEN out0_75 = to_unsigned(16#69#, 8) ELSE
      expandedKey(104);
  
  expandedKey_4(105) <= out0_105 WHEN out0_75 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(105);
  
  expandedKey_4(106) <= out0_105 WHEN out0_75 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(106);
  
  expandedKey_4(107) <= out0_105 WHEN out0_75 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(107);
  
  expandedKey_4(108) <= out0_105 WHEN out0_75 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(108);
  
  expandedKey_4(109) <= out0_105 WHEN out0_75 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(109);
  
  expandedKey_4(110) <= out0_105 WHEN out0_75 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(110);
  
  expandedKey_4(111) <= out0_105 WHEN out0_75 = to_unsigned(16#70#, 8) ELSE
      expandedKey(111);
  
  expandedKey_4(112) <= out0_105 WHEN out0_75 = to_unsigned(16#71#, 8) ELSE
      expandedKey(112);
  
  expandedKey_4(113) <= out0_105 WHEN out0_75 = to_unsigned(16#72#, 8) ELSE
      expandedKey(113);
  
  expandedKey_4(114) <= out0_105 WHEN out0_75 = to_unsigned(16#73#, 8) ELSE
      expandedKey(114);
  
  expandedKey_4(115) <= out0_105 WHEN out0_75 = to_unsigned(16#74#, 8) ELSE
      expandedKey(115);
  
  expandedKey_4(116) <= out0_105 WHEN out0_75 = to_unsigned(16#75#, 8) ELSE
      expandedKey(116);
  
  expandedKey_4(117) <= out0_105 WHEN out0_75 = to_unsigned(16#76#, 8) ELSE
      expandedKey(117);
  
  expandedKey_4(118) <= out0_105 WHEN out0_75 = to_unsigned(16#77#, 8) ELSE
      expandedKey(118);
  
  expandedKey_4(119) <= out0_105 WHEN out0_75 = to_unsigned(16#78#, 8) ELSE
      expandedKey(119);
  
  expandedKey_4(120) <= out0_105 WHEN out0_75 = to_unsigned(16#79#, 8) ELSE
      expandedKey(120);
  
  expandedKey_4(121) <= out0_105 WHEN out0_75 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(121);
  
  expandedKey_4(122) <= out0_105 WHEN out0_75 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(122);
  
  expandedKey_4(123) <= out0_105 WHEN out0_75 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(123);
  
  expandedKey_4(124) <= out0_105 WHEN out0_75 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(124);
  
  expandedKey_4(125) <= out0_105 WHEN out0_75 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(125);
  
  expandedKey_4(126) <= out0_105 WHEN out0_75 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(126);
  
  expandedKey_4(127) <= out0_105 WHEN out0_75 = to_unsigned(16#80#, 8) ELSE
      expandedKey(127);
  
  expandedKey_4(128) <= out0_105 WHEN out0_75 = to_unsigned(16#81#, 8) ELSE
      expandedKey(128);
  
  expandedKey_4(129) <= out0_105 WHEN out0_75 = to_unsigned(16#82#, 8) ELSE
      expandedKey(129);
  
  expandedKey_4(130) <= out0_105 WHEN out0_75 = to_unsigned(16#83#, 8) ELSE
      expandedKey(130);
  
  expandedKey_4(131) <= out0_105 WHEN out0_75 = to_unsigned(16#84#, 8) ELSE
      expandedKey(131);
  
  expandedKey_4(132) <= out0_105 WHEN out0_75 = to_unsigned(16#85#, 8) ELSE
      expandedKey(132);
  
  expandedKey_4(133) <= out0_105 WHEN out0_75 = to_unsigned(16#86#, 8) ELSE
      expandedKey(133);
  
  expandedKey_4(134) <= out0_105 WHEN out0_75 = to_unsigned(16#87#, 8) ELSE
      expandedKey(134);
  
  expandedKey_4(135) <= out0_105 WHEN out0_75 = to_unsigned(16#88#, 8) ELSE
      expandedKey(135);
  
  expandedKey_4(136) <= out0_105 WHEN out0_75 = to_unsigned(16#89#, 8) ELSE
      expandedKey(136);
  
  expandedKey_4(137) <= out0_105 WHEN out0_75 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(137);
  
  expandedKey_4(138) <= out0_105 WHEN out0_75 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(138);
  
  expandedKey_4(139) <= out0_105 WHEN out0_75 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(139);
  
  expandedKey_4(140) <= out0_105 WHEN out0_75 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(140);
  
  expandedKey_4(141) <= out0_105 WHEN out0_75 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(141);
  
  expandedKey_4(142) <= out0_105 WHEN out0_75 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(142);
  
  expandedKey_4(143) <= out0_105 WHEN out0_75 = to_unsigned(16#90#, 8) ELSE
      expandedKey(143);
  
  expandedKey_4(144) <= out0_105 WHEN out0_75 = to_unsigned(16#91#, 8) ELSE
      expandedKey(144);
  
  expandedKey_4(145) <= out0_105 WHEN out0_75 = to_unsigned(16#92#, 8) ELSE
      expandedKey(145);
  
  expandedKey_4(146) <= out0_105 WHEN out0_75 = to_unsigned(16#93#, 8) ELSE
      expandedKey(146);
  
  expandedKey_4(147) <= out0_105 WHEN out0_75 = to_unsigned(16#94#, 8) ELSE
      expandedKey(147);
  
  expandedKey_4(148) <= out0_105 WHEN out0_75 = to_unsigned(16#95#, 8) ELSE
      expandedKey(148);
  
  expandedKey_4(149) <= out0_105 WHEN out0_75 = to_unsigned(16#96#, 8) ELSE
      expandedKey(149);
  
  expandedKey_4(150) <= out0_105 WHEN out0_75 = to_unsigned(16#97#, 8) ELSE
      expandedKey(150);
  
  expandedKey_4(151) <= out0_105 WHEN out0_75 = to_unsigned(16#98#, 8) ELSE
      expandedKey(151);
  
  expandedKey_4(152) <= out0_105 WHEN out0_75 = to_unsigned(16#99#, 8) ELSE
      expandedKey(152);
  
  expandedKey_4(153) <= out0_105 WHEN out0_75 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(153);
  
  expandedKey_4(154) <= out0_105 WHEN out0_75 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(154);
  
  expandedKey_4(155) <= out0_105 WHEN out0_75 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(155);
  
  expandedKey_4(156) <= out0_105 WHEN out0_75 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(156);
  
  expandedKey_4(157) <= out0_105 WHEN out0_75 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(157);
  
  expandedKey_4(158) <= out0_105 WHEN out0_75 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(158);
  
  expandedKey_4(159) <= out0_105 WHEN out0_75 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(159);
  
  expandedKey_4(160) <= out0_105 WHEN out0_75 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(160);
  
  expandedKey_4(161) <= out0_105 WHEN out0_75 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(161);
  
  expandedKey_4(162) <= out0_105 WHEN out0_75 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(162);
  
  expandedKey_4(163) <= out0_105 WHEN out0_75 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(163);
  
  expandedKey_4(164) <= out0_105 WHEN out0_75 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(164);
  
  expandedKey_4(165) <= out0_105 WHEN out0_75 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(165);
  
  expandedKey_4(166) <= out0_105 WHEN out0_75 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(166);
  
  expandedKey_4(167) <= out0_105 WHEN out0_75 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(167);
  
  expandedKey_4(168) <= out0_105 WHEN out0_75 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(168);
  
  expandedKey_4(169) <= out0_105 WHEN out0_75 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(169);
  
  expandedKey_4(170) <= out0_105 WHEN out0_75 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(170);
  
  expandedKey_4(171) <= out0_105 WHEN out0_75 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(171);
  
  expandedKey_4(172) <= out0_105 WHEN out0_75 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(172);
  
  expandedKey_4(173) <= out0_105 WHEN out0_75 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(173);
  
  expandedKey_4(174) <= out0_105 WHEN out0_75 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(174);
  
  expandedKey_4(175) <= out0_105 WHEN out0_75 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(175);
  
  expandedKey_4(176) <= out0_105 WHEN out0_75 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(176);
  
  expandedKey_4(177) <= out0_105 WHEN out0_75 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(177);
  
  expandedKey_4(178) <= out0_105 WHEN out0_75 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(178);
  
  expandedKey_4(179) <= out0_105 WHEN out0_75 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(179);
  
  expandedKey_4(180) <= out0_105 WHEN out0_75 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(180);
  
  expandedKey_4(181) <= out0_105 WHEN out0_75 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(181);
  
  expandedKey_4(182) <= out0_105 WHEN out0_75 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(182);
  
  expandedKey_4(183) <= out0_105 WHEN out0_75 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(183);
  
  expandedKey_4(184) <= out0_105 WHEN out0_75 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(184);
  
  expandedKey_4(185) <= out0_105 WHEN out0_75 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(185);
  
  expandedKey_4(186) <= out0_105 WHEN out0_75 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(186);
  
  expandedKey_4(187) <= out0_105 WHEN out0_75 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(187);
  
  expandedKey_4(188) <= out0_105 WHEN out0_75 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(188);
  
  expandedKey_4(189) <= out0_105 WHEN out0_75 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(189);
  
  expandedKey_4(190) <= out0_105 WHEN out0_75 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(190);
  
  expandedKey_4(191) <= out0_105 WHEN out0_75 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(191);
  
  expandedKey_4(192) <= out0_105 WHEN out0_75 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(192);
  
  expandedKey_4(193) <= out0_105 WHEN out0_75 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(193);
  
  expandedKey_4(194) <= out0_105 WHEN out0_75 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(194);
  
  expandedKey_4(195) <= out0_105 WHEN out0_75 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(195);
  
  expandedKey_4(196) <= out0_105 WHEN out0_75 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(196);
  
  expandedKey_4(197) <= out0_105 WHEN out0_75 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(197);
  
  expandedKey_4(198) <= out0_105 WHEN out0_75 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(198);
  
  expandedKey_4(199) <= out0_105 WHEN out0_75 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(199);
  
  expandedKey_4(200) <= out0_105 WHEN out0_75 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(200);
  
  expandedKey_4(201) <= out0_105 WHEN out0_75 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(201);
  
  expandedKey_4(202) <= out0_105 WHEN out0_75 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(202);
  
  expandedKey_4(203) <= out0_105 WHEN out0_75 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(203);
  
  expandedKey_4(204) <= out0_105 WHEN out0_75 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(204);
  
  expandedKey_4(205) <= out0_105 WHEN out0_75 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(205);
  
  expandedKey_4(206) <= out0_105 WHEN out0_75 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(206);
  
  expandedKey_4(207) <= out0_105 WHEN out0_75 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(207);
  
  expandedKey_4(208) <= out0_105 WHEN out0_75 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(208);
  
  expandedKey_4(209) <= out0_105 WHEN out0_75 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(209);
  
  expandedKey_4(210) <= out0_105 WHEN out0_75 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(210);
  
  expandedKey_4(211) <= out0_105 WHEN out0_75 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(211);
  
  expandedKey_4(212) <= out0_105 WHEN out0_75 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(212);
  
  expandedKey_4(213) <= out0_105 WHEN out0_75 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(213);
  
  expandedKey_4(214) <= out0_105 WHEN out0_75 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(214);
  
  expandedKey_4(215) <= out0_105 WHEN out0_75 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(215);
  
  expandedKey_4(216) <= out0_105 WHEN out0_75 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(216);
  
  expandedKey_4(217) <= out0_105 WHEN out0_75 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(217);
  
  expandedKey_4(218) <= out0_105 WHEN out0_75 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(218);
  
  expandedKey_4(219) <= out0_105 WHEN out0_75 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(219);
  
  expandedKey_4(220) <= out0_105 WHEN out0_75 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(220);
  
  expandedKey_4(221) <= out0_105 WHEN out0_75 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(221);
  
  expandedKey_4(222) <= out0_105 WHEN out0_75 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(222);
  
  expandedKey_4(223) <= out0_105 WHEN out0_75 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(223);
  
  expandedKey_4(224) <= out0_105 WHEN out0_75 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(224);
  
  expandedKey_4(225) <= out0_105 WHEN out0_75 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(225);
  
  expandedKey_4(226) <= out0_105 WHEN out0_75 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(226);
  
  expandedKey_4(227) <= out0_105 WHEN out0_75 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(227);
  
  expandedKey_4(228) <= out0_105 WHEN out0_75 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(228);
  
  expandedKey_4(229) <= out0_105 WHEN out0_75 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(229);
  
  expandedKey_4(230) <= out0_105 WHEN out0_75 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(230);
  
  expandedKey_4(231) <= out0_105 WHEN out0_75 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(231);
  
  expandedKey_4(232) <= out0_105 WHEN out0_75 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(232);
  
  expandedKey_4(233) <= out0_105 WHEN out0_75 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(233);
  
  expandedKey_4(234) <= out0_105 WHEN out0_75 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(234);
  
  expandedKey_4(235) <= out0_105 WHEN out0_75 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(235);
  
  expandedKey_4(236) <= out0_105 WHEN out0_75 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(236);
  
  expandedKey_4(237) <= out0_105 WHEN out0_75 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(237);
  
  expandedKey_4(238) <= out0_105 WHEN out0_75 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(238);
  
  expandedKey_4(239) <= out0_105 WHEN out0_75 = to_unsigned(16#F0#, 8) ELSE
      expandedKey(239);

  
  expandedKey_3(0) <= out0_87 WHEN out0_77 = to_unsigned(16#01#, 8) ELSE
      expandedKey_4(0);
  
  expandedKey_3(1) <= out0_87 WHEN out0_77 = to_unsigned(16#02#, 8) ELSE
      expandedKey_4(1);
  
  expandedKey_3(2) <= out0_87 WHEN out0_77 = to_unsigned(16#03#, 8) ELSE
      expandedKey_4(2);
  
  expandedKey_3(3) <= out0_87 WHEN out0_77 = to_unsigned(16#04#, 8) ELSE
      expandedKey_4(3);
  
  expandedKey_3(4) <= out0_87 WHEN out0_77 = to_unsigned(16#05#, 8) ELSE
      expandedKey_4(4);
  
  expandedKey_3(5) <= out0_87 WHEN out0_77 = to_unsigned(16#06#, 8) ELSE
      expandedKey_4(5);
  
  expandedKey_3(6) <= out0_87 WHEN out0_77 = to_unsigned(16#07#, 8) ELSE
      expandedKey_4(6);
  
  expandedKey_3(7) <= out0_87 WHEN out0_77 = to_unsigned(16#08#, 8) ELSE
      expandedKey_4(7);
  
  expandedKey_3(8) <= out0_87 WHEN out0_77 = to_unsigned(16#09#, 8) ELSE
      expandedKey_4(8);
  
  expandedKey_3(9) <= out0_87 WHEN out0_77 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_4(9);
  
  expandedKey_3(10) <= out0_87 WHEN out0_77 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_4(10);
  
  expandedKey_3(11) <= out0_87 WHEN out0_77 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_4(11);
  
  expandedKey_3(12) <= out0_87 WHEN out0_77 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_4(12);
  
  expandedKey_3(13) <= out0_87 WHEN out0_77 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_4(13);
  
  expandedKey_3(14) <= out0_87 WHEN out0_77 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_4(14);
  
  expandedKey_3(15) <= out0_87 WHEN out0_77 = to_unsigned(16#10#, 8) ELSE
      expandedKey_4(15);
  
  expandedKey_3(16) <= out0_87 WHEN out0_77 = to_unsigned(16#11#, 8) ELSE
      expandedKey_4(16);
  
  expandedKey_3(17) <= out0_87 WHEN out0_77 = to_unsigned(16#12#, 8) ELSE
      expandedKey_4(17);
  
  expandedKey_3(18) <= out0_87 WHEN out0_77 = to_unsigned(16#13#, 8) ELSE
      expandedKey_4(18);
  
  expandedKey_3(19) <= out0_87 WHEN out0_77 = to_unsigned(16#14#, 8) ELSE
      expandedKey_4(19);
  
  expandedKey_3(20) <= out0_87 WHEN out0_77 = to_unsigned(16#15#, 8) ELSE
      expandedKey_4(20);
  
  expandedKey_3(21) <= out0_87 WHEN out0_77 = to_unsigned(16#16#, 8) ELSE
      expandedKey_4(21);
  
  expandedKey_3(22) <= out0_87 WHEN out0_77 = to_unsigned(16#17#, 8) ELSE
      expandedKey_4(22);
  
  expandedKey_3(23) <= out0_87 WHEN out0_77 = to_unsigned(16#18#, 8) ELSE
      expandedKey_4(23);
  
  expandedKey_3(24) <= out0_87 WHEN out0_77 = to_unsigned(16#19#, 8) ELSE
      expandedKey_4(24);
  
  expandedKey_3(25) <= out0_87 WHEN out0_77 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_4(25);
  
  expandedKey_3(26) <= out0_87 WHEN out0_77 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_4(26);
  
  expandedKey_3(27) <= out0_87 WHEN out0_77 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_4(27);
  
  expandedKey_3(28) <= out0_87 WHEN out0_77 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_4(28);
  
  expandedKey_3(29) <= out0_87 WHEN out0_77 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_4(29);
  
  expandedKey_3(30) <= out0_87 WHEN out0_77 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_4(30);
  
  expandedKey_3(31) <= out0_87 WHEN out0_77 = to_unsigned(16#20#, 8) ELSE
      expandedKey_4(31);
  
  expandedKey_3(32) <= out0_87 WHEN out0_77 = to_unsigned(16#21#, 8) ELSE
      expandedKey_4(32);
  
  expandedKey_3(33) <= out0_87 WHEN out0_77 = to_unsigned(16#22#, 8) ELSE
      expandedKey_4(33);
  
  expandedKey_3(34) <= out0_87 WHEN out0_77 = to_unsigned(16#23#, 8) ELSE
      expandedKey_4(34);
  
  expandedKey_3(35) <= out0_87 WHEN out0_77 = to_unsigned(16#24#, 8) ELSE
      expandedKey_4(35);
  
  expandedKey_3(36) <= out0_87 WHEN out0_77 = to_unsigned(16#25#, 8) ELSE
      expandedKey_4(36);
  
  expandedKey_3(37) <= out0_87 WHEN out0_77 = to_unsigned(16#26#, 8) ELSE
      expandedKey_4(37);
  
  expandedKey_3(38) <= out0_87 WHEN out0_77 = to_unsigned(16#27#, 8) ELSE
      expandedKey_4(38);
  
  expandedKey_3(39) <= out0_87 WHEN out0_77 = to_unsigned(16#28#, 8) ELSE
      expandedKey_4(39);
  
  expandedKey_3(40) <= out0_87 WHEN out0_77 = to_unsigned(16#29#, 8) ELSE
      expandedKey_4(40);
  
  expandedKey_3(41) <= out0_87 WHEN out0_77 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_4(41);
  
  expandedKey_3(42) <= out0_87 WHEN out0_77 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_4(42);
  
  expandedKey_3(43) <= out0_87 WHEN out0_77 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_4(43);
  
  expandedKey_3(44) <= out0_87 WHEN out0_77 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_4(44);
  
  expandedKey_3(45) <= out0_87 WHEN out0_77 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_4(45);
  
  expandedKey_3(46) <= out0_87 WHEN out0_77 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_4(46);
  
  expandedKey_3(47) <= out0_87 WHEN out0_77 = to_unsigned(16#30#, 8) ELSE
      expandedKey_4(47);
  
  expandedKey_3(48) <= out0_87 WHEN out0_77 = to_unsigned(16#31#, 8) ELSE
      expandedKey_4(48);
  
  expandedKey_3(49) <= out0_87 WHEN out0_77 = to_unsigned(16#32#, 8) ELSE
      expandedKey_4(49);
  
  expandedKey_3(50) <= out0_87 WHEN out0_77 = to_unsigned(16#33#, 8) ELSE
      expandedKey_4(50);
  
  expandedKey_3(51) <= out0_87 WHEN out0_77 = to_unsigned(16#34#, 8) ELSE
      expandedKey_4(51);
  
  expandedKey_3(52) <= out0_87 WHEN out0_77 = to_unsigned(16#35#, 8) ELSE
      expandedKey_4(52);
  
  expandedKey_3(53) <= out0_87 WHEN out0_77 = to_unsigned(16#36#, 8) ELSE
      expandedKey_4(53);
  
  expandedKey_3(54) <= out0_87 WHEN out0_77 = to_unsigned(16#37#, 8) ELSE
      expandedKey_4(54);
  
  expandedKey_3(55) <= out0_87 WHEN out0_77 = to_unsigned(16#38#, 8) ELSE
      expandedKey_4(55);
  
  expandedKey_3(56) <= out0_87 WHEN out0_77 = to_unsigned(16#39#, 8) ELSE
      expandedKey_4(56);
  
  expandedKey_3(57) <= out0_87 WHEN out0_77 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_4(57);
  
  expandedKey_3(58) <= out0_87 WHEN out0_77 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_4(58);
  
  expandedKey_3(59) <= out0_87 WHEN out0_77 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_4(59);
  
  expandedKey_3(60) <= out0_87 WHEN out0_77 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_4(60);
  
  expandedKey_3(61) <= out0_87 WHEN out0_77 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_4(61);
  
  expandedKey_3(62) <= out0_87 WHEN out0_77 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_4(62);
  
  expandedKey_3(63) <= out0_87 WHEN out0_77 = to_unsigned(16#40#, 8) ELSE
      expandedKey_4(63);
  
  expandedKey_3(64) <= out0_87 WHEN out0_77 = to_unsigned(16#41#, 8) ELSE
      expandedKey_4(64);
  
  expandedKey_3(65) <= out0_87 WHEN out0_77 = to_unsigned(16#42#, 8) ELSE
      expandedKey_4(65);
  
  expandedKey_3(66) <= out0_87 WHEN out0_77 = to_unsigned(16#43#, 8) ELSE
      expandedKey_4(66);
  
  expandedKey_3(67) <= out0_87 WHEN out0_77 = to_unsigned(16#44#, 8) ELSE
      expandedKey_4(67);
  
  expandedKey_3(68) <= out0_87 WHEN out0_77 = to_unsigned(16#45#, 8) ELSE
      expandedKey_4(68);
  
  expandedKey_3(69) <= out0_87 WHEN out0_77 = to_unsigned(16#46#, 8) ELSE
      expandedKey_4(69);
  
  expandedKey_3(70) <= out0_87 WHEN out0_77 = to_unsigned(16#47#, 8) ELSE
      expandedKey_4(70);
  
  expandedKey_3(71) <= out0_87 WHEN out0_77 = to_unsigned(16#48#, 8) ELSE
      expandedKey_4(71);
  
  expandedKey_3(72) <= out0_87 WHEN out0_77 = to_unsigned(16#49#, 8) ELSE
      expandedKey_4(72);
  
  expandedKey_3(73) <= out0_87 WHEN out0_77 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_4(73);
  
  expandedKey_3(74) <= out0_87 WHEN out0_77 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_4(74);
  
  expandedKey_3(75) <= out0_87 WHEN out0_77 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_4(75);
  
  expandedKey_3(76) <= out0_87 WHEN out0_77 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_4(76);
  
  expandedKey_3(77) <= out0_87 WHEN out0_77 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_4(77);
  
  expandedKey_3(78) <= out0_87 WHEN out0_77 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_4(78);
  
  expandedKey_3(79) <= out0_87 WHEN out0_77 = to_unsigned(16#50#, 8) ELSE
      expandedKey_4(79);
  
  expandedKey_3(80) <= out0_87 WHEN out0_77 = to_unsigned(16#51#, 8) ELSE
      expandedKey_4(80);
  
  expandedKey_3(81) <= out0_87 WHEN out0_77 = to_unsigned(16#52#, 8) ELSE
      expandedKey_4(81);
  
  expandedKey_3(82) <= out0_87 WHEN out0_77 = to_unsigned(16#53#, 8) ELSE
      expandedKey_4(82);
  
  expandedKey_3(83) <= out0_87 WHEN out0_77 = to_unsigned(16#54#, 8) ELSE
      expandedKey_4(83);
  
  expandedKey_3(84) <= out0_87 WHEN out0_77 = to_unsigned(16#55#, 8) ELSE
      expandedKey_4(84);
  
  expandedKey_3(85) <= out0_87 WHEN out0_77 = to_unsigned(16#56#, 8) ELSE
      expandedKey_4(85);
  
  expandedKey_3(86) <= out0_87 WHEN out0_77 = to_unsigned(16#57#, 8) ELSE
      expandedKey_4(86);
  
  expandedKey_3(87) <= out0_87 WHEN out0_77 = to_unsigned(16#58#, 8) ELSE
      expandedKey_4(87);
  
  expandedKey_3(88) <= out0_87 WHEN out0_77 = to_unsigned(16#59#, 8) ELSE
      expandedKey_4(88);
  
  expandedKey_3(89) <= out0_87 WHEN out0_77 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_4(89);
  
  expandedKey_3(90) <= out0_87 WHEN out0_77 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_4(90);
  
  expandedKey_3(91) <= out0_87 WHEN out0_77 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_4(91);
  
  expandedKey_3(92) <= out0_87 WHEN out0_77 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_4(92);
  
  expandedKey_3(93) <= out0_87 WHEN out0_77 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_4(93);
  
  expandedKey_3(94) <= out0_87 WHEN out0_77 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_4(94);
  
  expandedKey_3(95) <= out0_87 WHEN out0_77 = to_unsigned(16#60#, 8) ELSE
      expandedKey_4(95);
  
  expandedKey_3(96) <= out0_87 WHEN out0_77 = to_unsigned(16#61#, 8) ELSE
      expandedKey_4(96);
  
  expandedKey_3(97) <= out0_87 WHEN out0_77 = to_unsigned(16#62#, 8) ELSE
      expandedKey_4(97);
  
  expandedKey_3(98) <= out0_87 WHEN out0_77 = to_unsigned(16#63#, 8) ELSE
      expandedKey_4(98);
  
  expandedKey_3(99) <= out0_87 WHEN out0_77 = to_unsigned(16#64#, 8) ELSE
      expandedKey_4(99);
  
  expandedKey_3(100) <= out0_87 WHEN out0_77 = to_unsigned(16#65#, 8) ELSE
      expandedKey_4(100);
  
  expandedKey_3(101) <= out0_87 WHEN out0_77 = to_unsigned(16#66#, 8) ELSE
      expandedKey_4(101);
  
  expandedKey_3(102) <= out0_87 WHEN out0_77 = to_unsigned(16#67#, 8) ELSE
      expandedKey_4(102);
  
  expandedKey_3(103) <= out0_87 WHEN out0_77 = to_unsigned(16#68#, 8) ELSE
      expandedKey_4(103);
  
  expandedKey_3(104) <= out0_87 WHEN out0_77 = to_unsigned(16#69#, 8) ELSE
      expandedKey_4(104);
  
  expandedKey_3(105) <= out0_87 WHEN out0_77 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_4(105);
  
  expandedKey_3(106) <= out0_87 WHEN out0_77 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_4(106);
  
  expandedKey_3(107) <= out0_87 WHEN out0_77 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_4(107);
  
  expandedKey_3(108) <= out0_87 WHEN out0_77 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_4(108);
  
  expandedKey_3(109) <= out0_87 WHEN out0_77 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_4(109);
  
  expandedKey_3(110) <= out0_87 WHEN out0_77 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_4(110);
  
  expandedKey_3(111) <= out0_87 WHEN out0_77 = to_unsigned(16#70#, 8) ELSE
      expandedKey_4(111);
  
  expandedKey_3(112) <= out0_87 WHEN out0_77 = to_unsigned(16#71#, 8) ELSE
      expandedKey_4(112);
  
  expandedKey_3(113) <= out0_87 WHEN out0_77 = to_unsigned(16#72#, 8) ELSE
      expandedKey_4(113);
  
  expandedKey_3(114) <= out0_87 WHEN out0_77 = to_unsigned(16#73#, 8) ELSE
      expandedKey_4(114);
  
  expandedKey_3(115) <= out0_87 WHEN out0_77 = to_unsigned(16#74#, 8) ELSE
      expandedKey_4(115);
  
  expandedKey_3(116) <= out0_87 WHEN out0_77 = to_unsigned(16#75#, 8) ELSE
      expandedKey_4(116);
  
  expandedKey_3(117) <= out0_87 WHEN out0_77 = to_unsigned(16#76#, 8) ELSE
      expandedKey_4(117);
  
  expandedKey_3(118) <= out0_87 WHEN out0_77 = to_unsigned(16#77#, 8) ELSE
      expandedKey_4(118);
  
  expandedKey_3(119) <= out0_87 WHEN out0_77 = to_unsigned(16#78#, 8) ELSE
      expandedKey_4(119);
  
  expandedKey_3(120) <= out0_87 WHEN out0_77 = to_unsigned(16#79#, 8) ELSE
      expandedKey_4(120);
  
  expandedKey_3(121) <= out0_87 WHEN out0_77 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_4(121);
  
  expandedKey_3(122) <= out0_87 WHEN out0_77 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_4(122);
  
  expandedKey_3(123) <= out0_87 WHEN out0_77 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_4(123);
  
  expandedKey_3(124) <= out0_87 WHEN out0_77 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_4(124);
  
  expandedKey_3(125) <= out0_87 WHEN out0_77 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_4(125);
  
  expandedKey_3(126) <= out0_87 WHEN out0_77 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_4(126);
  
  expandedKey_3(127) <= out0_87 WHEN out0_77 = to_unsigned(16#80#, 8) ELSE
      expandedKey_4(127);
  
  expandedKey_3(128) <= out0_87 WHEN out0_77 = to_unsigned(16#81#, 8) ELSE
      expandedKey_4(128);
  
  expandedKey_3(129) <= out0_87 WHEN out0_77 = to_unsigned(16#82#, 8) ELSE
      expandedKey_4(129);
  
  expandedKey_3(130) <= out0_87 WHEN out0_77 = to_unsigned(16#83#, 8) ELSE
      expandedKey_4(130);
  
  expandedKey_3(131) <= out0_87 WHEN out0_77 = to_unsigned(16#84#, 8) ELSE
      expandedKey_4(131);
  
  expandedKey_3(132) <= out0_87 WHEN out0_77 = to_unsigned(16#85#, 8) ELSE
      expandedKey_4(132);
  
  expandedKey_3(133) <= out0_87 WHEN out0_77 = to_unsigned(16#86#, 8) ELSE
      expandedKey_4(133);
  
  expandedKey_3(134) <= out0_87 WHEN out0_77 = to_unsigned(16#87#, 8) ELSE
      expandedKey_4(134);
  
  expandedKey_3(135) <= out0_87 WHEN out0_77 = to_unsigned(16#88#, 8) ELSE
      expandedKey_4(135);
  
  expandedKey_3(136) <= out0_87 WHEN out0_77 = to_unsigned(16#89#, 8) ELSE
      expandedKey_4(136);
  
  expandedKey_3(137) <= out0_87 WHEN out0_77 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_4(137);
  
  expandedKey_3(138) <= out0_87 WHEN out0_77 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_4(138);
  
  expandedKey_3(139) <= out0_87 WHEN out0_77 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_4(139);
  
  expandedKey_3(140) <= out0_87 WHEN out0_77 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_4(140);
  
  expandedKey_3(141) <= out0_87 WHEN out0_77 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_4(141);
  
  expandedKey_3(142) <= out0_87 WHEN out0_77 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_4(142);
  
  expandedKey_3(143) <= out0_87 WHEN out0_77 = to_unsigned(16#90#, 8) ELSE
      expandedKey_4(143);
  
  expandedKey_3(144) <= out0_87 WHEN out0_77 = to_unsigned(16#91#, 8) ELSE
      expandedKey_4(144);
  
  expandedKey_3(145) <= out0_87 WHEN out0_77 = to_unsigned(16#92#, 8) ELSE
      expandedKey_4(145);
  
  expandedKey_3(146) <= out0_87 WHEN out0_77 = to_unsigned(16#93#, 8) ELSE
      expandedKey_4(146);
  
  expandedKey_3(147) <= out0_87 WHEN out0_77 = to_unsigned(16#94#, 8) ELSE
      expandedKey_4(147);
  
  expandedKey_3(148) <= out0_87 WHEN out0_77 = to_unsigned(16#95#, 8) ELSE
      expandedKey_4(148);
  
  expandedKey_3(149) <= out0_87 WHEN out0_77 = to_unsigned(16#96#, 8) ELSE
      expandedKey_4(149);
  
  expandedKey_3(150) <= out0_87 WHEN out0_77 = to_unsigned(16#97#, 8) ELSE
      expandedKey_4(150);
  
  expandedKey_3(151) <= out0_87 WHEN out0_77 = to_unsigned(16#98#, 8) ELSE
      expandedKey_4(151);
  
  expandedKey_3(152) <= out0_87 WHEN out0_77 = to_unsigned(16#99#, 8) ELSE
      expandedKey_4(152);
  
  expandedKey_3(153) <= out0_87 WHEN out0_77 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_4(153);
  
  expandedKey_3(154) <= out0_87 WHEN out0_77 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_4(154);
  
  expandedKey_3(155) <= out0_87 WHEN out0_77 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_4(155);
  
  expandedKey_3(156) <= out0_87 WHEN out0_77 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_4(156);
  
  expandedKey_3(157) <= out0_87 WHEN out0_77 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_4(157);
  
  expandedKey_3(158) <= out0_87 WHEN out0_77 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_4(158);
  
  expandedKey_3(159) <= out0_87 WHEN out0_77 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_4(159);
  
  expandedKey_3(160) <= out0_87 WHEN out0_77 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_4(160);
  
  expandedKey_3(161) <= out0_87 WHEN out0_77 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_4(161);
  
  expandedKey_3(162) <= out0_87 WHEN out0_77 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_4(162);
  
  expandedKey_3(163) <= out0_87 WHEN out0_77 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_4(163);
  
  expandedKey_3(164) <= out0_87 WHEN out0_77 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_4(164);
  
  expandedKey_3(165) <= out0_87 WHEN out0_77 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_4(165);
  
  expandedKey_3(166) <= out0_87 WHEN out0_77 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_4(166);
  
  expandedKey_3(167) <= out0_87 WHEN out0_77 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_4(167);
  
  expandedKey_3(168) <= out0_87 WHEN out0_77 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_4(168);
  
  expandedKey_3(169) <= out0_87 WHEN out0_77 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_4(169);
  
  expandedKey_3(170) <= out0_87 WHEN out0_77 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_4(170);
  
  expandedKey_3(171) <= out0_87 WHEN out0_77 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_4(171);
  
  expandedKey_3(172) <= out0_87 WHEN out0_77 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_4(172);
  
  expandedKey_3(173) <= out0_87 WHEN out0_77 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_4(173);
  
  expandedKey_3(174) <= out0_87 WHEN out0_77 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_4(174);
  
  expandedKey_3(175) <= out0_87 WHEN out0_77 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_4(175);
  
  expandedKey_3(176) <= out0_87 WHEN out0_77 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_4(176);
  
  expandedKey_3(177) <= out0_87 WHEN out0_77 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_4(177);
  
  expandedKey_3(178) <= out0_87 WHEN out0_77 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_4(178);
  
  expandedKey_3(179) <= out0_87 WHEN out0_77 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_4(179);
  
  expandedKey_3(180) <= out0_87 WHEN out0_77 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_4(180);
  
  expandedKey_3(181) <= out0_87 WHEN out0_77 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_4(181);
  
  expandedKey_3(182) <= out0_87 WHEN out0_77 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_4(182);
  
  expandedKey_3(183) <= out0_87 WHEN out0_77 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_4(183);
  
  expandedKey_3(184) <= out0_87 WHEN out0_77 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_4(184);
  
  expandedKey_3(185) <= out0_87 WHEN out0_77 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_4(185);
  
  expandedKey_3(186) <= out0_87 WHEN out0_77 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_4(186);
  
  expandedKey_3(187) <= out0_87 WHEN out0_77 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_4(187);
  
  expandedKey_3(188) <= out0_87 WHEN out0_77 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_4(188);
  
  expandedKey_3(189) <= out0_87 WHEN out0_77 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_4(189);
  
  expandedKey_3(190) <= out0_87 WHEN out0_77 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_4(190);
  
  expandedKey_3(191) <= out0_87 WHEN out0_77 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_4(191);
  
  expandedKey_3(192) <= out0_87 WHEN out0_77 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_4(192);
  
  expandedKey_3(193) <= out0_87 WHEN out0_77 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_4(193);
  
  expandedKey_3(194) <= out0_87 WHEN out0_77 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_4(194);
  
  expandedKey_3(195) <= out0_87 WHEN out0_77 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_4(195);
  
  expandedKey_3(196) <= out0_87 WHEN out0_77 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_4(196);
  
  expandedKey_3(197) <= out0_87 WHEN out0_77 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_4(197);
  
  expandedKey_3(198) <= out0_87 WHEN out0_77 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_4(198);
  
  expandedKey_3(199) <= out0_87 WHEN out0_77 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_4(199);
  
  expandedKey_3(200) <= out0_87 WHEN out0_77 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_4(200);
  
  expandedKey_3(201) <= out0_87 WHEN out0_77 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_4(201);
  
  expandedKey_3(202) <= out0_87 WHEN out0_77 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_4(202);
  
  expandedKey_3(203) <= out0_87 WHEN out0_77 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_4(203);
  
  expandedKey_3(204) <= out0_87 WHEN out0_77 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_4(204);
  
  expandedKey_3(205) <= out0_87 WHEN out0_77 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_4(205);
  
  expandedKey_3(206) <= out0_87 WHEN out0_77 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_4(206);
  
  expandedKey_3(207) <= out0_87 WHEN out0_77 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_4(207);
  
  expandedKey_3(208) <= out0_87 WHEN out0_77 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_4(208);
  
  expandedKey_3(209) <= out0_87 WHEN out0_77 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_4(209);
  
  expandedKey_3(210) <= out0_87 WHEN out0_77 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_4(210);
  
  expandedKey_3(211) <= out0_87 WHEN out0_77 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_4(211);
  
  expandedKey_3(212) <= out0_87 WHEN out0_77 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_4(212);
  
  expandedKey_3(213) <= out0_87 WHEN out0_77 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_4(213);
  
  expandedKey_3(214) <= out0_87 WHEN out0_77 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_4(214);
  
  expandedKey_3(215) <= out0_87 WHEN out0_77 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_4(215);
  
  expandedKey_3(216) <= out0_87 WHEN out0_77 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_4(216);
  
  expandedKey_3(217) <= out0_87 WHEN out0_77 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_4(217);
  
  expandedKey_3(218) <= out0_87 WHEN out0_77 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_4(218);
  
  expandedKey_3(219) <= out0_87 WHEN out0_77 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_4(219);
  
  expandedKey_3(220) <= out0_87 WHEN out0_77 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_4(220);
  
  expandedKey_3(221) <= out0_87 WHEN out0_77 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_4(221);
  
  expandedKey_3(222) <= out0_87 WHEN out0_77 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_4(222);
  
  expandedKey_3(223) <= out0_87 WHEN out0_77 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_4(223);
  
  expandedKey_3(224) <= out0_87 WHEN out0_77 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_4(224);
  
  expandedKey_3(225) <= out0_87 WHEN out0_77 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_4(225);
  
  expandedKey_3(226) <= out0_87 WHEN out0_77 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_4(226);
  
  expandedKey_3(227) <= out0_87 WHEN out0_77 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_4(227);
  
  expandedKey_3(228) <= out0_87 WHEN out0_77 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_4(228);
  
  expandedKey_3(229) <= out0_87 WHEN out0_77 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_4(229);
  
  expandedKey_3(230) <= out0_87 WHEN out0_77 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_4(230);
  
  expandedKey_3(231) <= out0_87 WHEN out0_77 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_4(231);
  
  expandedKey_3(232) <= out0_87 WHEN out0_77 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_4(232);
  
  expandedKey_3(233) <= out0_87 WHEN out0_77 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_4(233);
  
  expandedKey_3(234) <= out0_87 WHEN out0_77 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_4(234);
  
  expandedKey_3(235) <= out0_87 WHEN out0_77 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_4(235);
  
  expandedKey_3(236) <= out0_87 WHEN out0_77 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_4(236);
  
  expandedKey_3(237) <= out0_87 WHEN out0_77 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_4(237);
  
  expandedKey_3(238) <= out0_87 WHEN out0_77 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_4(238);
  
  expandedKey_3(239) <= out0_87 WHEN out0_77 = to_unsigned(16#F0#, 8) ELSE
      expandedKey_4(239);

  
  expandedKey_2(0) <= out0_85 WHEN out0_79 = to_unsigned(16#01#, 8) ELSE
      expandedKey_3(0);
  
  expandedKey_2(1) <= out0_85 WHEN out0_79 = to_unsigned(16#02#, 8) ELSE
      expandedKey_3(1);
  
  expandedKey_2(2) <= out0_85 WHEN out0_79 = to_unsigned(16#03#, 8) ELSE
      expandedKey_3(2);
  
  expandedKey_2(3) <= out0_85 WHEN out0_79 = to_unsigned(16#04#, 8) ELSE
      expandedKey_3(3);
  
  expandedKey_2(4) <= out0_85 WHEN out0_79 = to_unsigned(16#05#, 8) ELSE
      expandedKey_3(4);
  
  expandedKey_2(5) <= out0_85 WHEN out0_79 = to_unsigned(16#06#, 8) ELSE
      expandedKey_3(5);
  
  expandedKey_2(6) <= out0_85 WHEN out0_79 = to_unsigned(16#07#, 8) ELSE
      expandedKey_3(6);
  
  expandedKey_2(7) <= out0_85 WHEN out0_79 = to_unsigned(16#08#, 8) ELSE
      expandedKey_3(7);
  
  expandedKey_2(8) <= out0_85 WHEN out0_79 = to_unsigned(16#09#, 8) ELSE
      expandedKey_3(8);
  
  expandedKey_2(9) <= out0_85 WHEN out0_79 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_3(9);
  
  expandedKey_2(10) <= out0_85 WHEN out0_79 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_3(10);
  
  expandedKey_2(11) <= out0_85 WHEN out0_79 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_3(11);
  
  expandedKey_2(12) <= out0_85 WHEN out0_79 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_3(12);
  
  expandedKey_2(13) <= out0_85 WHEN out0_79 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_3(13);
  
  expandedKey_2(14) <= out0_85 WHEN out0_79 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_3(14);
  
  expandedKey_2(15) <= out0_85 WHEN out0_79 = to_unsigned(16#10#, 8) ELSE
      expandedKey_3(15);
  
  expandedKey_2(16) <= out0_85 WHEN out0_79 = to_unsigned(16#11#, 8) ELSE
      expandedKey_3(16);
  
  expandedKey_2(17) <= out0_85 WHEN out0_79 = to_unsigned(16#12#, 8) ELSE
      expandedKey_3(17);
  
  expandedKey_2(18) <= out0_85 WHEN out0_79 = to_unsigned(16#13#, 8) ELSE
      expandedKey_3(18);
  
  expandedKey_2(19) <= out0_85 WHEN out0_79 = to_unsigned(16#14#, 8) ELSE
      expandedKey_3(19);
  
  expandedKey_2(20) <= out0_85 WHEN out0_79 = to_unsigned(16#15#, 8) ELSE
      expandedKey_3(20);
  
  expandedKey_2(21) <= out0_85 WHEN out0_79 = to_unsigned(16#16#, 8) ELSE
      expandedKey_3(21);
  
  expandedKey_2(22) <= out0_85 WHEN out0_79 = to_unsigned(16#17#, 8) ELSE
      expandedKey_3(22);
  
  expandedKey_2(23) <= out0_85 WHEN out0_79 = to_unsigned(16#18#, 8) ELSE
      expandedKey_3(23);
  
  expandedKey_2(24) <= out0_85 WHEN out0_79 = to_unsigned(16#19#, 8) ELSE
      expandedKey_3(24);
  
  expandedKey_2(25) <= out0_85 WHEN out0_79 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_3(25);
  
  expandedKey_2(26) <= out0_85 WHEN out0_79 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_3(26);
  
  expandedKey_2(27) <= out0_85 WHEN out0_79 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_3(27);
  
  expandedKey_2(28) <= out0_85 WHEN out0_79 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_3(28);
  
  expandedKey_2(29) <= out0_85 WHEN out0_79 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_3(29);
  
  expandedKey_2(30) <= out0_85 WHEN out0_79 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_3(30);
  
  expandedKey_2(31) <= out0_85 WHEN out0_79 = to_unsigned(16#20#, 8) ELSE
      expandedKey_3(31);
  
  expandedKey_2(32) <= out0_85 WHEN out0_79 = to_unsigned(16#21#, 8) ELSE
      expandedKey_3(32);
  
  expandedKey_2(33) <= out0_85 WHEN out0_79 = to_unsigned(16#22#, 8) ELSE
      expandedKey_3(33);
  
  expandedKey_2(34) <= out0_85 WHEN out0_79 = to_unsigned(16#23#, 8) ELSE
      expandedKey_3(34);
  
  expandedKey_2(35) <= out0_85 WHEN out0_79 = to_unsigned(16#24#, 8) ELSE
      expandedKey_3(35);
  
  expandedKey_2(36) <= out0_85 WHEN out0_79 = to_unsigned(16#25#, 8) ELSE
      expandedKey_3(36);
  
  expandedKey_2(37) <= out0_85 WHEN out0_79 = to_unsigned(16#26#, 8) ELSE
      expandedKey_3(37);
  
  expandedKey_2(38) <= out0_85 WHEN out0_79 = to_unsigned(16#27#, 8) ELSE
      expandedKey_3(38);
  
  expandedKey_2(39) <= out0_85 WHEN out0_79 = to_unsigned(16#28#, 8) ELSE
      expandedKey_3(39);
  
  expandedKey_2(40) <= out0_85 WHEN out0_79 = to_unsigned(16#29#, 8) ELSE
      expandedKey_3(40);
  
  expandedKey_2(41) <= out0_85 WHEN out0_79 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_3(41);
  
  expandedKey_2(42) <= out0_85 WHEN out0_79 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_3(42);
  
  expandedKey_2(43) <= out0_85 WHEN out0_79 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_3(43);
  
  expandedKey_2(44) <= out0_85 WHEN out0_79 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_3(44);
  
  expandedKey_2(45) <= out0_85 WHEN out0_79 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_3(45);
  
  expandedKey_2(46) <= out0_85 WHEN out0_79 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_3(46);
  
  expandedKey_2(47) <= out0_85 WHEN out0_79 = to_unsigned(16#30#, 8) ELSE
      expandedKey_3(47);
  
  expandedKey_2(48) <= out0_85 WHEN out0_79 = to_unsigned(16#31#, 8) ELSE
      expandedKey_3(48);
  
  expandedKey_2(49) <= out0_85 WHEN out0_79 = to_unsigned(16#32#, 8) ELSE
      expandedKey_3(49);
  
  expandedKey_2(50) <= out0_85 WHEN out0_79 = to_unsigned(16#33#, 8) ELSE
      expandedKey_3(50);
  
  expandedKey_2(51) <= out0_85 WHEN out0_79 = to_unsigned(16#34#, 8) ELSE
      expandedKey_3(51);
  
  expandedKey_2(52) <= out0_85 WHEN out0_79 = to_unsigned(16#35#, 8) ELSE
      expandedKey_3(52);
  
  expandedKey_2(53) <= out0_85 WHEN out0_79 = to_unsigned(16#36#, 8) ELSE
      expandedKey_3(53);
  
  expandedKey_2(54) <= out0_85 WHEN out0_79 = to_unsigned(16#37#, 8) ELSE
      expandedKey_3(54);
  
  expandedKey_2(55) <= out0_85 WHEN out0_79 = to_unsigned(16#38#, 8) ELSE
      expandedKey_3(55);
  
  expandedKey_2(56) <= out0_85 WHEN out0_79 = to_unsigned(16#39#, 8) ELSE
      expandedKey_3(56);
  
  expandedKey_2(57) <= out0_85 WHEN out0_79 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_3(57);
  
  expandedKey_2(58) <= out0_85 WHEN out0_79 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_3(58);
  
  expandedKey_2(59) <= out0_85 WHEN out0_79 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_3(59);
  
  expandedKey_2(60) <= out0_85 WHEN out0_79 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_3(60);
  
  expandedKey_2(61) <= out0_85 WHEN out0_79 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_3(61);
  
  expandedKey_2(62) <= out0_85 WHEN out0_79 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_3(62);
  
  expandedKey_2(63) <= out0_85 WHEN out0_79 = to_unsigned(16#40#, 8) ELSE
      expandedKey_3(63);
  
  expandedKey_2(64) <= out0_85 WHEN out0_79 = to_unsigned(16#41#, 8) ELSE
      expandedKey_3(64);
  
  expandedKey_2(65) <= out0_85 WHEN out0_79 = to_unsigned(16#42#, 8) ELSE
      expandedKey_3(65);
  
  expandedKey_2(66) <= out0_85 WHEN out0_79 = to_unsigned(16#43#, 8) ELSE
      expandedKey_3(66);
  
  expandedKey_2(67) <= out0_85 WHEN out0_79 = to_unsigned(16#44#, 8) ELSE
      expandedKey_3(67);
  
  expandedKey_2(68) <= out0_85 WHEN out0_79 = to_unsigned(16#45#, 8) ELSE
      expandedKey_3(68);
  
  expandedKey_2(69) <= out0_85 WHEN out0_79 = to_unsigned(16#46#, 8) ELSE
      expandedKey_3(69);
  
  expandedKey_2(70) <= out0_85 WHEN out0_79 = to_unsigned(16#47#, 8) ELSE
      expandedKey_3(70);
  
  expandedKey_2(71) <= out0_85 WHEN out0_79 = to_unsigned(16#48#, 8) ELSE
      expandedKey_3(71);
  
  expandedKey_2(72) <= out0_85 WHEN out0_79 = to_unsigned(16#49#, 8) ELSE
      expandedKey_3(72);
  
  expandedKey_2(73) <= out0_85 WHEN out0_79 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_3(73);
  
  expandedKey_2(74) <= out0_85 WHEN out0_79 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_3(74);
  
  expandedKey_2(75) <= out0_85 WHEN out0_79 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_3(75);
  
  expandedKey_2(76) <= out0_85 WHEN out0_79 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_3(76);
  
  expandedKey_2(77) <= out0_85 WHEN out0_79 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_3(77);
  
  expandedKey_2(78) <= out0_85 WHEN out0_79 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_3(78);
  
  expandedKey_2(79) <= out0_85 WHEN out0_79 = to_unsigned(16#50#, 8) ELSE
      expandedKey_3(79);
  
  expandedKey_2(80) <= out0_85 WHEN out0_79 = to_unsigned(16#51#, 8) ELSE
      expandedKey_3(80);
  
  expandedKey_2(81) <= out0_85 WHEN out0_79 = to_unsigned(16#52#, 8) ELSE
      expandedKey_3(81);
  
  expandedKey_2(82) <= out0_85 WHEN out0_79 = to_unsigned(16#53#, 8) ELSE
      expandedKey_3(82);
  
  expandedKey_2(83) <= out0_85 WHEN out0_79 = to_unsigned(16#54#, 8) ELSE
      expandedKey_3(83);
  
  expandedKey_2(84) <= out0_85 WHEN out0_79 = to_unsigned(16#55#, 8) ELSE
      expandedKey_3(84);
  
  expandedKey_2(85) <= out0_85 WHEN out0_79 = to_unsigned(16#56#, 8) ELSE
      expandedKey_3(85);
  
  expandedKey_2(86) <= out0_85 WHEN out0_79 = to_unsigned(16#57#, 8) ELSE
      expandedKey_3(86);
  
  expandedKey_2(87) <= out0_85 WHEN out0_79 = to_unsigned(16#58#, 8) ELSE
      expandedKey_3(87);
  
  expandedKey_2(88) <= out0_85 WHEN out0_79 = to_unsigned(16#59#, 8) ELSE
      expandedKey_3(88);
  
  expandedKey_2(89) <= out0_85 WHEN out0_79 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_3(89);
  
  expandedKey_2(90) <= out0_85 WHEN out0_79 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_3(90);
  
  expandedKey_2(91) <= out0_85 WHEN out0_79 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_3(91);
  
  expandedKey_2(92) <= out0_85 WHEN out0_79 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_3(92);
  
  expandedKey_2(93) <= out0_85 WHEN out0_79 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_3(93);
  
  expandedKey_2(94) <= out0_85 WHEN out0_79 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_3(94);
  
  expandedKey_2(95) <= out0_85 WHEN out0_79 = to_unsigned(16#60#, 8) ELSE
      expandedKey_3(95);
  
  expandedKey_2(96) <= out0_85 WHEN out0_79 = to_unsigned(16#61#, 8) ELSE
      expandedKey_3(96);
  
  expandedKey_2(97) <= out0_85 WHEN out0_79 = to_unsigned(16#62#, 8) ELSE
      expandedKey_3(97);
  
  expandedKey_2(98) <= out0_85 WHEN out0_79 = to_unsigned(16#63#, 8) ELSE
      expandedKey_3(98);
  
  expandedKey_2(99) <= out0_85 WHEN out0_79 = to_unsigned(16#64#, 8) ELSE
      expandedKey_3(99);
  
  expandedKey_2(100) <= out0_85 WHEN out0_79 = to_unsigned(16#65#, 8) ELSE
      expandedKey_3(100);
  
  expandedKey_2(101) <= out0_85 WHEN out0_79 = to_unsigned(16#66#, 8) ELSE
      expandedKey_3(101);
  
  expandedKey_2(102) <= out0_85 WHEN out0_79 = to_unsigned(16#67#, 8) ELSE
      expandedKey_3(102);
  
  expandedKey_2(103) <= out0_85 WHEN out0_79 = to_unsigned(16#68#, 8) ELSE
      expandedKey_3(103);
  
  expandedKey_2(104) <= out0_85 WHEN out0_79 = to_unsigned(16#69#, 8) ELSE
      expandedKey_3(104);
  
  expandedKey_2(105) <= out0_85 WHEN out0_79 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_3(105);
  
  expandedKey_2(106) <= out0_85 WHEN out0_79 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_3(106);
  
  expandedKey_2(107) <= out0_85 WHEN out0_79 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_3(107);
  
  expandedKey_2(108) <= out0_85 WHEN out0_79 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_3(108);
  
  expandedKey_2(109) <= out0_85 WHEN out0_79 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_3(109);
  
  expandedKey_2(110) <= out0_85 WHEN out0_79 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_3(110);
  
  expandedKey_2(111) <= out0_85 WHEN out0_79 = to_unsigned(16#70#, 8) ELSE
      expandedKey_3(111);
  
  expandedKey_2(112) <= out0_85 WHEN out0_79 = to_unsigned(16#71#, 8) ELSE
      expandedKey_3(112);
  
  expandedKey_2(113) <= out0_85 WHEN out0_79 = to_unsigned(16#72#, 8) ELSE
      expandedKey_3(113);
  
  expandedKey_2(114) <= out0_85 WHEN out0_79 = to_unsigned(16#73#, 8) ELSE
      expandedKey_3(114);
  
  expandedKey_2(115) <= out0_85 WHEN out0_79 = to_unsigned(16#74#, 8) ELSE
      expandedKey_3(115);
  
  expandedKey_2(116) <= out0_85 WHEN out0_79 = to_unsigned(16#75#, 8) ELSE
      expandedKey_3(116);
  
  expandedKey_2(117) <= out0_85 WHEN out0_79 = to_unsigned(16#76#, 8) ELSE
      expandedKey_3(117);
  
  expandedKey_2(118) <= out0_85 WHEN out0_79 = to_unsigned(16#77#, 8) ELSE
      expandedKey_3(118);
  
  expandedKey_2(119) <= out0_85 WHEN out0_79 = to_unsigned(16#78#, 8) ELSE
      expandedKey_3(119);
  
  expandedKey_2(120) <= out0_85 WHEN out0_79 = to_unsigned(16#79#, 8) ELSE
      expandedKey_3(120);
  
  expandedKey_2(121) <= out0_85 WHEN out0_79 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_3(121);
  
  expandedKey_2(122) <= out0_85 WHEN out0_79 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_3(122);
  
  expandedKey_2(123) <= out0_85 WHEN out0_79 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_3(123);
  
  expandedKey_2(124) <= out0_85 WHEN out0_79 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_3(124);
  
  expandedKey_2(125) <= out0_85 WHEN out0_79 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_3(125);
  
  expandedKey_2(126) <= out0_85 WHEN out0_79 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_3(126);
  
  expandedKey_2(127) <= out0_85 WHEN out0_79 = to_unsigned(16#80#, 8) ELSE
      expandedKey_3(127);
  
  expandedKey_2(128) <= out0_85 WHEN out0_79 = to_unsigned(16#81#, 8) ELSE
      expandedKey_3(128);
  
  expandedKey_2(129) <= out0_85 WHEN out0_79 = to_unsigned(16#82#, 8) ELSE
      expandedKey_3(129);
  
  expandedKey_2(130) <= out0_85 WHEN out0_79 = to_unsigned(16#83#, 8) ELSE
      expandedKey_3(130);
  
  expandedKey_2(131) <= out0_85 WHEN out0_79 = to_unsigned(16#84#, 8) ELSE
      expandedKey_3(131);
  
  expandedKey_2(132) <= out0_85 WHEN out0_79 = to_unsigned(16#85#, 8) ELSE
      expandedKey_3(132);
  
  expandedKey_2(133) <= out0_85 WHEN out0_79 = to_unsigned(16#86#, 8) ELSE
      expandedKey_3(133);
  
  expandedKey_2(134) <= out0_85 WHEN out0_79 = to_unsigned(16#87#, 8) ELSE
      expandedKey_3(134);
  
  expandedKey_2(135) <= out0_85 WHEN out0_79 = to_unsigned(16#88#, 8) ELSE
      expandedKey_3(135);
  
  expandedKey_2(136) <= out0_85 WHEN out0_79 = to_unsigned(16#89#, 8) ELSE
      expandedKey_3(136);
  
  expandedKey_2(137) <= out0_85 WHEN out0_79 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_3(137);
  
  expandedKey_2(138) <= out0_85 WHEN out0_79 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_3(138);
  
  expandedKey_2(139) <= out0_85 WHEN out0_79 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_3(139);
  
  expandedKey_2(140) <= out0_85 WHEN out0_79 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_3(140);
  
  expandedKey_2(141) <= out0_85 WHEN out0_79 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_3(141);
  
  expandedKey_2(142) <= out0_85 WHEN out0_79 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_3(142);
  
  expandedKey_2(143) <= out0_85 WHEN out0_79 = to_unsigned(16#90#, 8) ELSE
      expandedKey_3(143);
  
  expandedKey_2(144) <= out0_85 WHEN out0_79 = to_unsigned(16#91#, 8) ELSE
      expandedKey_3(144);
  
  expandedKey_2(145) <= out0_85 WHEN out0_79 = to_unsigned(16#92#, 8) ELSE
      expandedKey_3(145);
  
  expandedKey_2(146) <= out0_85 WHEN out0_79 = to_unsigned(16#93#, 8) ELSE
      expandedKey_3(146);
  
  expandedKey_2(147) <= out0_85 WHEN out0_79 = to_unsigned(16#94#, 8) ELSE
      expandedKey_3(147);
  
  expandedKey_2(148) <= out0_85 WHEN out0_79 = to_unsigned(16#95#, 8) ELSE
      expandedKey_3(148);
  
  expandedKey_2(149) <= out0_85 WHEN out0_79 = to_unsigned(16#96#, 8) ELSE
      expandedKey_3(149);
  
  expandedKey_2(150) <= out0_85 WHEN out0_79 = to_unsigned(16#97#, 8) ELSE
      expandedKey_3(150);
  
  expandedKey_2(151) <= out0_85 WHEN out0_79 = to_unsigned(16#98#, 8) ELSE
      expandedKey_3(151);
  
  expandedKey_2(152) <= out0_85 WHEN out0_79 = to_unsigned(16#99#, 8) ELSE
      expandedKey_3(152);
  
  expandedKey_2(153) <= out0_85 WHEN out0_79 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_3(153);
  
  expandedKey_2(154) <= out0_85 WHEN out0_79 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_3(154);
  
  expandedKey_2(155) <= out0_85 WHEN out0_79 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_3(155);
  
  expandedKey_2(156) <= out0_85 WHEN out0_79 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_3(156);
  
  expandedKey_2(157) <= out0_85 WHEN out0_79 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_3(157);
  
  expandedKey_2(158) <= out0_85 WHEN out0_79 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_3(158);
  
  expandedKey_2(159) <= out0_85 WHEN out0_79 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_3(159);
  
  expandedKey_2(160) <= out0_85 WHEN out0_79 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_3(160);
  
  expandedKey_2(161) <= out0_85 WHEN out0_79 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_3(161);
  
  expandedKey_2(162) <= out0_85 WHEN out0_79 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_3(162);
  
  expandedKey_2(163) <= out0_85 WHEN out0_79 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_3(163);
  
  expandedKey_2(164) <= out0_85 WHEN out0_79 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_3(164);
  
  expandedKey_2(165) <= out0_85 WHEN out0_79 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_3(165);
  
  expandedKey_2(166) <= out0_85 WHEN out0_79 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_3(166);
  
  expandedKey_2(167) <= out0_85 WHEN out0_79 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_3(167);
  
  expandedKey_2(168) <= out0_85 WHEN out0_79 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_3(168);
  
  expandedKey_2(169) <= out0_85 WHEN out0_79 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_3(169);
  
  expandedKey_2(170) <= out0_85 WHEN out0_79 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_3(170);
  
  expandedKey_2(171) <= out0_85 WHEN out0_79 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_3(171);
  
  expandedKey_2(172) <= out0_85 WHEN out0_79 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_3(172);
  
  expandedKey_2(173) <= out0_85 WHEN out0_79 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_3(173);
  
  expandedKey_2(174) <= out0_85 WHEN out0_79 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_3(174);
  
  expandedKey_2(175) <= out0_85 WHEN out0_79 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_3(175);
  
  expandedKey_2(176) <= out0_85 WHEN out0_79 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_3(176);
  
  expandedKey_2(177) <= out0_85 WHEN out0_79 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_3(177);
  
  expandedKey_2(178) <= out0_85 WHEN out0_79 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_3(178);
  
  expandedKey_2(179) <= out0_85 WHEN out0_79 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_3(179);
  
  expandedKey_2(180) <= out0_85 WHEN out0_79 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_3(180);
  
  expandedKey_2(181) <= out0_85 WHEN out0_79 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_3(181);
  
  expandedKey_2(182) <= out0_85 WHEN out0_79 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_3(182);
  
  expandedKey_2(183) <= out0_85 WHEN out0_79 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_3(183);
  
  expandedKey_2(184) <= out0_85 WHEN out0_79 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_3(184);
  
  expandedKey_2(185) <= out0_85 WHEN out0_79 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_3(185);
  
  expandedKey_2(186) <= out0_85 WHEN out0_79 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_3(186);
  
  expandedKey_2(187) <= out0_85 WHEN out0_79 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_3(187);
  
  expandedKey_2(188) <= out0_85 WHEN out0_79 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_3(188);
  
  expandedKey_2(189) <= out0_85 WHEN out0_79 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_3(189);
  
  expandedKey_2(190) <= out0_85 WHEN out0_79 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_3(190);
  
  expandedKey_2(191) <= out0_85 WHEN out0_79 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_3(191);
  
  expandedKey_2(192) <= out0_85 WHEN out0_79 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_3(192);
  
  expandedKey_2(193) <= out0_85 WHEN out0_79 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_3(193);
  
  expandedKey_2(194) <= out0_85 WHEN out0_79 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_3(194);
  
  expandedKey_2(195) <= out0_85 WHEN out0_79 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_3(195);
  
  expandedKey_2(196) <= out0_85 WHEN out0_79 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_3(196);
  
  expandedKey_2(197) <= out0_85 WHEN out0_79 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_3(197);
  
  expandedKey_2(198) <= out0_85 WHEN out0_79 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_3(198);
  
  expandedKey_2(199) <= out0_85 WHEN out0_79 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_3(199);
  
  expandedKey_2(200) <= out0_85 WHEN out0_79 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_3(200);
  
  expandedKey_2(201) <= out0_85 WHEN out0_79 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_3(201);
  
  expandedKey_2(202) <= out0_85 WHEN out0_79 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_3(202);
  
  expandedKey_2(203) <= out0_85 WHEN out0_79 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_3(203);
  
  expandedKey_2(204) <= out0_85 WHEN out0_79 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_3(204);
  
  expandedKey_2(205) <= out0_85 WHEN out0_79 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_3(205);
  
  expandedKey_2(206) <= out0_85 WHEN out0_79 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_3(206);
  
  expandedKey_2(207) <= out0_85 WHEN out0_79 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_3(207);
  
  expandedKey_2(208) <= out0_85 WHEN out0_79 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_3(208);
  
  expandedKey_2(209) <= out0_85 WHEN out0_79 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_3(209);
  
  expandedKey_2(210) <= out0_85 WHEN out0_79 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_3(210);
  
  expandedKey_2(211) <= out0_85 WHEN out0_79 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_3(211);
  
  expandedKey_2(212) <= out0_85 WHEN out0_79 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_3(212);
  
  expandedKey_2(213) <= out0_85 WHEN out0_79 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_3(213);
  
  expandedKey_2(214) <= out0_85 WHEN out0_79 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_3(214);
  
  expandedKey_2(215) <= out0_85 WHEN out0_79 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_3(215);
  
  expandedKey_2(216) <= out0_85 WHEN out0_79 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_3(216);
  
  expandedKey_2(217) <= out0_85 WHEN out0_79 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_3(217);
  
  expandedKey_2(218) <= out0_85 WHEN out0_79 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_3(218);
  
  expandedKey_2(219) <= out0_85 WHEN out0_79 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_3(219);
  
  expandedKey_2(220) <= out0_85 WHEN out0_79 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_3(220);
  
  expandedKey_2(221) <= out0_85 WHEN out0_79 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_3(221);
  
  expandedKey_2(222) <= out0_85 WHEN out0_79 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_3(222);
  
  expandedKey_2(223) <= out0_85 WHEN out0_79 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_3(223);
  
  expandedKey_2(224) <= out0_85 WHEN out0_79 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_3(224);
  
  expandedKey_2(225) <= out0_85 WHEN out0_79 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_3(225);
  
  expandedKey_2(226) <= out0_85 WHEN out0_79 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_3(226);
  
  expandedKey_2(227) <= out0_85 WHEN out0_79 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_3(227);
  
  expandedKey_2(228) <= out0_85 WHEN out0_79 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_3(228);
  
  expandedKey_2(229) <= out0_85 WHEN out0_79 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_3(229);
  
  expandedKey_2(230) <= out0_85 WHEN out0_79 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_3(230);
  
  expandedKey_2(231) <= out0_85 WHEN out0_79 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_3(231);
  
  expandedKey_2(232) <= out0_85 WHEN out0_79 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_3(232);
  
  expandedKey_2(233) <= out0_85 WHEN out0_79 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_3(233);
  
  expandedKey_2(234) <= out0_85 WHEN out0_79 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_3(234);
  
  expandedKey_2(235) <= out0_85 WHEN out0_79 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_3(235);
  
  expandedKey_2(236) <= out0_85 WHEN out0_79 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_3(236);
  
  expandedKey_2(237) <= out0_85 WHEN out0_79 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_3(237);
  
  expandedKey_2(238) <= out0_85 WHEN out0_79 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_3(238);
  
  expandedKey_2(239) <= out0_85 WHEN out0_79 = to_unsigned(16#F0#, 8) ELSE
      expandedKey_3(239);

  
  expandedKey_5(0) <= out0_83 WHEN out0_81 = to_unsigned(16#01#, 8) ELSE
      expandedKey_2(0);
  
  expandedKey_5(1) <= out0_83 WHEN out0_81 = to_unsigned(16#02#, 8) ELSE
      expandedKey_2(1);
  
  expandedKey_5(2) <= out0_83 WHEN out0_81 = to_unsigned(16#03#, 8) ELSE
      expandedKey_2(2);
  
  expandedKey_5(3) <= out0_83 WHEN out0_81 = to_unsigned(16#04#, 8) ELSE
      expandedKey_2(3);
  
  expandedKey_5(4) <= out0_83 WHEN out0_81 = to_unsigned(16#05#, 8) ELSE
      expandedKey_2(4);
  
  expandedKey_5(5) <= out0_83 WHEN out0_81 = to_unsigned(16#06#, 8) ELSE
      expandedKey_2(5);
  
  expandedKey_5(6) <= out0_83 WHEN out0_81 = to_unsigned(16#07#, 8) ELSE
      expandedKey_2(6);
  
  expandedKey_5(7) <= out0_83 WHEN out0_81 = to_unsigned(16#08#, 8) ELSE
      expandedKey_2(7);
  
  expandedKey_5(8) <= out0_83 WHEN out0_81 = to_unsigned(16#09#, 8) ELSE
      expandedKey_2(8);
  
  expandedKey_5(9) <= out0_83 WHEN out0_81 = to_unsigned(16#0A#, 8) ELSE
      expandedKey_2(9);
  
  expandedKey_5(10) <= out0_83 WHEN out0_81 = to_unsigned(16#0B#, 8) ELSE
      expandedKey_2(10);
  
  expandedKey_5(11) <= out0_83 WHEN out0_81 = to_unsigned(16#0C#, 8) ELSE
      expandedKey_2(11);
  
  expandedKey_5(12) <= out0_83 WHEN out0_81 = to_unsigned(16#0D#, 8) ELSE
      expandedKey_2(12);
  
  expandedKey_5(13) <= out0_83 WHEN out0_81 = to_unsigned(16#0E#, 8) ELSE
      expandedKey_2(13);
  
  expandedKey_5(14) <= out0_83 WHEN out0_81 = to_unsigned(16#0F#, 8) ELSE
      expandedKey_2(14);
  
  expandedKey_5(15) <= out0_83 WHEN out0_81 = to_unsigned(16#10#, 8) ELSE
      expandedKey_2(15);
  
  expandedKey_5(16) <= out0_83 WHEN out0_81 = to_unsigned(16#11#, 8) ELSE
      expandedKey_2(16);
  
  expandedKey_5(17) <= out0_83 WHEN out0_81 = to_unsigned(16#12#, 8) ELSE
      expandedKey_2(17);
  
  expandedKey_5(18) <= out0_83 WHEN out0_81 = to_unsigned(16#13#, 8) ELSE
      expandedKey_2(18);
  
  expandedKey_5(19) <= out0_83 WHEN out0_81 = to_unsigned(16#14#, 8) ELSE
      expandedKey_2(19);
  
  expandedKey_5(20) <= out0_83 WHEN out0_81 = to_unsigned(16#15#, 8) ELSE
      expandedKey_2(20);
  
  expandedKey_5(21) <= out0_83 WHEN out0_81 = to_unsigned(16#16#, 8) ELSE
      expandedKey_2(21);
  
  expandedKey_5(22) <= out0_83 WHEN out0_81 = to_unsigned(16#17#, 8) ELSE
      expandedKey_2(22);
  
  expandedKey_5(23) <= out0_83 WHEN out0_81 = to_unsigned(16#18#, 8) ELSE
      expandedKey_2(23);
  
  expandedKey_5(24) <= out0_83 WHEN out0_81 = to_unsigned(16#19#, 8) ELSE
      expandedKey_2(24);
  
  expandedKey_5(25) <= out0_83 WHEN out0_81 = to_unsigned(16#1A#, 8) ELSE
      expandedKey_2(25);
  
  expandedKey_5(26) <= out0_83 WHEN out0_81 = to_unsigned(16#1B#, 8) ELSE
      expandedKey_2(26);
  
  expandedKey_5(27) <= out0_83 WHEN out0_81 = to_unsigned(16#1C#, 8) ELSE
      expandedKey_2(27);
  
  expandedKey_5(28) <= out0_83 WHEN out0_81 = to_unsigned(16#1D#, 8) ELSE
      expandedKey_2(28);
  
  expandedKey_5(29) <= out0_83 WHEN out0_81 = to_unsigned(16#1E#, 8) ELSE
      expandedKey_2(29);
  
  expandedKey_5(30) <= out0_83 WHEN out0_81 = to_unsigned(16#1F#, 8) ELSE
      expandedKey_2(30);
  
  expandedKey_5(31) <= out0_83 WHEN out0_81 = to_unsigned(16#20#, 8) ELSE
      expandedKey_2(31);
  
  expandedKey_5(32) <= out0_83 WHEN out0_81 = to_unsigned(16#21#, 8) ELSE
      expandedKey_2(32);
  
  expandedKey_5(33) <= out0_83 WHEN out0_81 = to_unsigned(16#22#, 8) ELSE
      expandedKey_2(33);
  
  expandedKey_5(34) <= out0_83 WHEN out0_81 = to_unsigned(16#23#, 8) ELSE
      expandedKey_2(34);
  
  expandedKey_5(35) <= out0_83 WHEN out0_81 = to_unsigned(16#24#, 8) ELSE
      expandedKey_2(35);
  
  expandedKey_5(36) <= out0_83 WHEN out0_81 = to_unsigned(16#25#, 8) ELSE
      expandedKey_2(36);
  
  expandedKey_5(37) <= out0_83 WHEN out0_81 = to_unsigned(16#26#, 8) ELSE
      expandedKey_2(37);
  
  expandedKey_5(38) <= out0_83 WHEN out0_81 = to_unsigned(16#27#, 8) ELSE
      expandedKey_2(38);
  
  expandedKey_5(39) <= out0_83 WHEN out0_81 = to_unsigned(16#28#, 8) ELSE
      expandedKey_2(39);
  
  expandedKey_5(40) <= out0_83 WHEN out0_81 = to_unsigned(16#29#, 8) ELSE
      expandedKey_2(40);
  
  expandedKey_5(41) <= out0_83 WHEN out0_81 = to_unsigned(16#2A#, 8) ELSE
      expandedKey_2(41);
  
  expandedKey_5(42) <= out0_83 WHEN out0_81 = to_unsigned(16#2B#, 8) ELSE
      expandedKey_2(42);
  
  expandedKey_5(43) <= out0_83 WHEN out0_81 = to_unsigned(16#2C#, 8) ELSE
      expandedKey_2(43);
  
  expandedKey_5(44) <= out0_83 WHEN out0_81 = to_unsigned(16#2D#, 8) ELSE
      expandedKey_2(44);
  
  expandedKey_5(45) <= out0_83 WHEN out0_81 = to_unsigned(16#2E#, 8) ELSE
      expandedKey_2(45);
  
  expandedKey_5(46) <= out0_83 WHEN out0_81 = to_unsigned(16#2F#, 8) ELSE
      expandedKey_2(46);
  
  expandedKey_5(47) <= out0_83 WHEN out0_81 = to_unsigned(16#30#, 8) ELSE
      expandedKey_2(47);
  
  expandedKey_5(48) <= out0_83 WHEN out0_81 = to_unsigned(16#31#, 8) ELSE
      expandedKey_2(48);
  
  expandedKey_5(49) <= out0_83 WHEN out0_81 = to_unsigned(16#32#, 8) ELSE
      expandedKey_2(49);
  
  expandedKey_5(50) <= out0_83 WHEN out0_81 = to_unsigned(16#33#, 8) ELSE
      expandedKey_2(50);
  
  expandedKey_5(51) <= out0_83 WHEN out0_81 = to_unsigned(16#34#, 8) ELSE
      expandedKey_2(51);
  
  expandedKey_5(52) <= out0_83 WHEN out0_81 = to_unsigned(16#35#, 8) ELSE
      expandedKey_2(52);
  
  expandedKey_5(53) <= out0_83 WHEN out0_81 = to_unsigned(16#36#, 8) ELSE
      expandedKey_2(53);
  
  expandedKey_5(54) <= out0_83 WHEN out0_81 = to_unsigned(16#37#, 8) ELSE
      expandedKey_2(54);
  
  expandedKey_5(55) <= out0_83 WHEN out0_81 = to_unsigned(16#38#, 8) ELSE
      expandedKey_2(55);
  
  expandedKey_5(56) <= out0_83 WHEN out0_81 = to_unsigned(16#39#, 8) ELSE
      expandedKey_2(56);
  
  expandedKey_5(57) <= out0_83 WHEN out0_81 = to_unsigned(16#3A#, 8) ELSE
      expandedKey_2(57);
  
  expandedKey_5(58) <= out0_83 WHEN out0_81 = to_unsigned(16#3B#, 8) ELSE
      expandedKey_2(58);
  
  expandedKey_5(59) <= out0_83 WHEN out0_81 = to_unsigned(16#3C#, 8) ELSE
      expandedKey_2(59);
  
  expandedKey_5(60) <= out0_83 WHEN out0_81 = to_unsigned(16#3D#, 8) ELSE
      expandedKey_2(60);
  
  expandedKey_5(61) <= out0_83 WHEN out0_81 = to_unsigned(16#3E#, 8) ELSE
      expandedKey_2(61);
  
  expandedKey_5(62) <= out0_83 WHEN out0_81 = to_unsigned(16#3F#, 8) ELSE
      expandedKey_2(62);
  
  expandedKey_5(63) <= out0_83 WHEN out0_81 = to_unsigned(16#40#, 8) ELSE
      expandedKey_2(63);
  
  expandedKey_5(64) <= out0_83 WHEN out0_81 = to_unsigned(16#41#, 8) ELSE
      expandedKey_2(64);
  
  expandedKey_5(65) <= out0_83 WHEN out0_81 = to_unsigned(16#42#, 8) ELSE
      expandedKey_2(65);
  
  expandedKey_5(66) <= out0_83 WHEN out0_81 = to_unsigned(16#43#, 8) ELSE
      expandedKey_2(66);
  
  expandedKey_5(67) <= out0_83 WHEN out0_81 = to_unsigned(16#44#, 8) ELSE
      expandedKey_2(67);
  
  expandedKey_5(68) <= out0_83 WHEN out0_81 = to_unsigned(16#45#, 8) ELSE
      expandedKey_2(68);
  
  expandedKey_5(69) <= out0_83 WHEN out0_81 = to_unsigned(16#46#, 8) ELSE
      expandedKey_2(69);
  
  expandedKey_5(70) <= out0_83 WHEN out0_81 = to_unsigned(16#47#, 8) ELSE
      expandedKey_2(70);
  
  expandedKey_5(71) <= out0_83 WHEN out0_81 = to_unsigned(16#48#, 8) ELSE
      expandedKey_2(71);
  
  expandedKey_5(72) <= out0_83 WHEN out0_81 = to_unsigned(16#49#, 8) ELSE
      expandedKey_2(72);
  
  expandedKey_5(73) <= out0_83 WHEN out0_81 = to_unsigned(16#4A#, 8) ELSE
      expandedKey_2(73);
  
  expandedKey_5(74) <= out0_83 WHEN out0_81 = to_unsigned(16#4B#, 8) ELSE
      expandedKey_2(74);
  
  expandedKey_5(75) <= out0_83 WHEN out0_81 = to_unsigned(16#4C#, 8) ELSE
      expandedKey_2(75);
  
  expandedKey_5(76) <= out0_83 WHEN out0_81 = to_unsigned(16#4D#, 8) ELSE
      expandedKey_2(76);
  
  expandedKey_5(77) <= out0_83 WHEN out0_81 = to_unsigned(16#4E#, 8) ELSE
      expandedKey_2(77);
  
  expandedKey_5(78) <= out0_83 WHEN out0_81 = to_unsigned(16#4F#, 8) ELSE
      expandedKey_2(78);
  
  expandedKey_5(79) <= out0_83 WHEN out0_81 = to_unsigned(16#50#, 8) ELSE
      expandedKey_2(79);
  
  expandedKey_5(80) <= out0_83 WHEN out0_81 = to_unsigned(16#51#, 8) ELSE
      expandedKey_2(80);
  
  expandedKey_5(81) <= out0_83 WHEN out0_81 = to_unsigned(16#52#, 8) ELSE
      expandedKey_2(81);
  
  expandedKey_5(82) <= out0_83 WHEN out0_81 = to_unsigned(16#53#, 8) ELSE
      expandedKey_2(82);
  
  expandedKey_5(83) <= out0_83 WHEN out0_81 = to_unsigned(16#54#, 8) ELSE
      expandedKey_2(83);
  
  expandedKey_5(84) <= out0_83 WHEN out0_81 = to_unsigned(16#55#, 8) ELSE
      expandedKey_2(84);
  
  expandedKey_5(85) <= out0_83 WHEN out0_81 = to_unsigned(16#56#, 8) ELSE
      expandedKey_2(85);
  
  expandedKey_5(86) <= out0_83 WHEN out0_81 = to_unsigned(16#57#, 8) ELSE
      expandedKey_2(86);
  
  expandedKey_5(87) <= out0_83 WHEN out0_81 = to_unsigned(16#58#, 8) ELSE
      expandedKey_2(87);
  
  expandedKey_5(88) <= out0_83 WHEN out0_81 = to_unsigned(16#59#, 8) ELSE
      expandedKey_2(88);
  
  expandedKey_5(89) <= out0_83 WHEN out0_81 = to_unsigned(16#5A#, 8) ELSE
      expandedKey_2(89);
  
  expandedKey_5(90) <= out0_83 WHEN out0_81 = to_unsigned(16#5B#, 8) ELSE
      expandedKey_2(90);
  
  expandedKey_5(91) <= out0_83 WHEN out0_81 = to_unsigned(16#5C#, 8) ELSE
      expandedKey_2(91);
  
  expandedKey_5(92) <= out0_83 WHEN out0_81 = to_unsigned(16#5D#, 8) ELSE
      expandedKey_2(92);
  
  expandedKey_5(93) <= out0_83 WHEN out0_81 = to_unsigned(16#5E#, 8) ELSE
      expandedKey_2(93);
  
  expandedKey_5(94) <= out0_83 WHEN out0_81 = to_unsigned(16#5F#, 8) ELSE
      expandedKey_2(94);
  
  expandedKey_5(95) <= out0_83 WHEN out0_81 = to_unsigned(16#60#, 8) ELSE
      expandedKey_2(95);
  
  expandedKey_5(96) <= out0_83 WHEN out0_81 = to_unsigned(16#61#, 8) ELSE
      expandedKey_2(96);
  
  expandedKey_5(97) <= out0_83 WHEN out0_81 = to_unsigned(16#62#, 8) ELSE
      expandedKey_2(97);
  
  expandedKey_5(98) <= out0_83 WHEN out0_81 = to_unsigned(16#63#, 8) ELSE
      expandedKey_2(98);
  
  expandedKey_5(99) <= out0_83 WHEN out0_81 = to_unsigned(16#64#, 8) ELSE
      expandedKey_2(99);
  
  expandedKey_5(100) <= out0_83 WHEN out0_81 = to_unsigned(16#65#, 8) ELSE
      expandedKey_2(100);
  
  expandedKey_5(101) <= out0_83 WHEN out0_81 = to_unsigned(16#66#, 8) ELSE
      expandedKey_2(101);
  
  expandedKey_5(102) <= out0_83 WHEN out0_81 = to_unsigned(16#67#, 8) ELSE
      expandedKey_2(102);
  
  expandedKey_5(103) <= out0_83 WHEN out0_81 = to_unsigned(16#68#, 8) ELSE
      expandedKey_2(103);
  
  expandedKey_5(104) <= out0_83 WHEN out0_81 = to_unsigned(16#69#, 8) ELSE
      expandedKey_2(104);
  
  expandedKey_5(105) <= out0_83 WHEN out0_81 = to_unsigned(16#6A#, 8) ELSE
      expandedKey_2(105);
  
  expandedKey_5(106) <= out0_83 WHEN out0_81 = to_unsigned(16#6B#, 8) ELSE
      expandedKey_2(106);
  
  expandedKey_5(107) <= out0_83 WHEN out0_81 = to_unsigned(16#6C#, 8) ELSE
      expandedKey_2(107);
  
  expandedKey_5(108) <= out0_83 WHEN out0_81 = to_unsigned(16#6D#, 8) ELSE
      expandedKey_2(108);
  
  expandedKey_5(109) <= out0_83 WHEN out0_81 = to_unsigned(16#6E#, 8) ELSE
      expandedKey_2(109);
  
  expandedKey_5(110) <= out0_83 WHEN out0_81 = to_unsigned(16#6F#, 8) ELSE
      expandedKey_2(110);
  
  expandedKey_5(111) <= out0_83 WHEN out0_81 = to_unsigned(16#70#, 8) ELSE
      expandedKey_2(111);
  
  expandedKey_5(112) <= out0_83 WHEN out0_81 = to_unsigned(16#71#, 8) ELSE
      expandedKey_2(112);
  
  expandedKey_5(113) <= out0_83 WHEN out0_81 = to_unsigned(16#72#, 8) ELSE
      expandedKey_2(113);
  
  expandedKey_5(114) <= out0_83 WHEN out0_81 = to_unsigned(16#73#, 8) ELSE
      expandedKey_2(114);
  
  expandedKey_5(115) <= out0_83 WHEN out0_81 = to_unsigned(16#74#, 8) ELSE
      expandedKey_2(115);
  
  expandedKey_5(116) <= out0_83 WHEN out0_81 = to_unsigned(16#75#, 8) ELSE
      expandedKey_2(116);
  
  expandedKey_5(117) <= out0_83 WHEN out0_81 = to_unsigned(16#76#, 8) ELSE
      expandedKey_2(117);
  
  expandedKey_5(118) <= out0_83 WHEN out0_81 = to_unsigned(16#77#, 8) ELSE
      expandedKey_2(118);
  
  expandedKey_5(119) <= out0_83 WHEN out0_81 = to_unsigned(16#78#, 8) ELSE
      expandedKey_2(119);
  
  expandedKey_5(120) <= out0_83 WHEN out0_81 = to_unsigned(16#79#, 8) ELSE
      expandedKey_2(120);
  
  expandedKey_5(121) <= out0_83 WHEN out0_81 = to_unsigned(16#7A#, 8) ELSE
      expandedKey_2(121);
  
  expandedKey_5(122) <= out0_83 WHEN out0_81 = to_unsigned(16#7B#, 8) ELSE
      expandedKey_2(122);
  
  expandedKey_5(123) <= out0_83 WHEN out0_81 = to_unsigned(16#7C#, 8) ELSE
      expandedKey_2(123);
  
  expandedKey_5(124) <= out0_83 WHEN out0_81 = to_unsigned(16#7D#, 8) ELSE
      expandedKey_2(124);
  
  expandedKey_5(125) <= out0_83 WHEN out0_81 = to_unsigned(16#7E#, 8) ELSE
      expandedKey_2(125);
  
  expandedKey_5(126) <= out0_83 WHEN out0_81 = to_unsigned(16#7F#, 8) ELSE
      expandedKey_2(126);
  
  expandedKey_5(127) <= out0_83 WHEN out0_81 = to_unsigned(16#80#, 8) ELSE
      expandedKey_2(127);
  
  expandedKey_5(128) <= out0_83 WHEN out0_81 = to_unsigned(16#81#, 8) ELSE
      expandedKey_2(128);
  
  expandedKey_5(129) <= out0_83 WHEN out0_81 = to_unsigned(16#82#, 8) ELSE
      expandedKey_2(129);
  
  expandedKey_5(130) <= out0_83 WHEN out0_81 = to_unsigned(16#83#, 8) ELSE
      expandedKey_2(130);
  
  expandedKey_5(131) <= out0_83 WHEN out0_81 = to_unsigned(16#84#, 8) ELSE
      expandedKey_2(131);
  
  expandedKey_5(132) <= out0_83 WHEN out0_81 = to_unsigned(16#85#, 8) ELSE
      expandedKey_2(132);
  
  expandedKey_5(133) <= out0_83 WHEN out0_81 = to_unsigned(16#86#, 8) ELSE
      expandedKey_2(133);
  
  expandedKey_5(134) <= out0_83 WHEN out0_81 = to_unsigned(16#87#, 8) ELSE
      expandedKey_2(134);
  
  expandedKey_5(135) <= out0_83 WHEN out0_81 = to_unsigned(16#88#, 8) ELSE
      expandedKey_2(135);
  
  expandedKey_5(136) <= out0_83 WHEN out0_81 = to_unsigned(16#89#, 8) ELSE
      expandedKey_2(136);
  
  expandedKey_5(137) <= out0_83 WHEN out0_81 = to_unsigned(16#8A#, 8) ELSE
      expandedKey_2(137);
  
  expandedKey_5(138) <= out0_83 WHEN out0_81 = to_unsigned(16#8B#, 8) ELSE
      expandedKey_2(138);
  
  expandedKey_5(139) <= out0_83 WHEN out0_81 = to_unsigned(16#8C#, 8) ELSE
      expandedKey_2(139);
  
  expandedKey_5(140) <= out0_83 WHEN out0_81 = to_unsigned(16#8D#, 8) ELSE
      expandedKey_2(140);
  
  expandedKey_5(141) <= out0_83 WHEN out0_81 = to_unsigned(16#8E#, 8) ELSE
      expandedKey_2(141);
  
  expandedKey_5(142) <= out0_83 WHEN out0_81 = to_unsigned(16#8F#, 8) ELSE
      expandedKey_2(142);
  
  expandedKey_5(143) <= out0_83 WHEN out0_81 = to_unsigned(16#90#, 8) ELSE
      expandedKey_2(143);
  
  expandedKey_5(144) <= out0_83 WHEN out0_81 = to_unsigned(16#91#, 8) ELSE
      expandedKey_2(144);
  
  expandedKey_5(145) <= out0_83 WHEN out0_81 = to_unsigned(16#92#, 8) ELSE
      expandedKey_2(145);
  
  expandedKey_5(146) <= out0_83 WHEN out0_81 = to_unsigned(16#93#, 8) ELSE
      expandedKey_2(146);
  
  expandedKey_5(147) <= out0_83 WHEN out0_81 = to_unsigned(16#94#, 8) ELSE
      expandedKey_2(147);
  
  expandedKey_5(148) <= out0_83 WHEN out0_81 = to_unsigned(16#95#, 8) ELSE
      expandedKey_2(148);
  
  expandedKey_5(149) <= out0_83 WHEN out0_81 = to_unsigned(16#96#, 8) ELSE
      expandedKey_2(149);
  
  expandedKey_5(150) <= out0_83 WHEN out0_81 = to_unsigned(16#97#, 8) ELSE
      expandedKey_2(150);
  
  expandedKey_5(151) <= out0_83 WHEN out0_81 = to_unsigned(16#98#, 8) ELSE
      expandedKey_2(151);
  
  expandedKey_5(152) <= out0_83 WHEN out0_81 = to_unsigned(16#99#, 8) ELSE
      expandedKey_2(152);
  
  expandedKey_5(153) <= out0_83 WHEN out0_81 = to_unsigned(16#9A#, 8) ELSE
      expandedKey_2(153);
  
  expandedKey_5(154) <= out0_83 WHEN out0_81 = to_unsigned(16#9B#, 8) ELSE
      expandedKey_2(154);
  
  expandedKey_5(155) <= out0_83 WHEN out0_81 = to_unsigned(16#9C#, 8) ELSE
      expandedKey_2(155);
  
  expandedKey_5(156) <= out0_83 WHEN out0_81 = to_unsigned(16#9D#, 8) ELSE
      expandedKey_2(156);
  
  expandedKey_5(157) <= out0_83 WHEN out0_81 = to_unsigned(16#9E#, 8) ELSE
      expandedKey_2(157);
  
  expandedKey_5(158) <= out0_83 WHEN out0_81 = to_unsigned(16#9F#, 8) ELSE
      expandedKey_2(158);
  
  expandedKey_5(159) <= out0_83 WHEN out0_81 = to_unsigned(16#A0#, 8) ELSE
      expandedKey_2(159);
  
  expandedKey_5(160) <= out0_83 WHEN out0_81 = to_unsigned(16#A1#, 8) ELSE
      expandedKey_2(160);
  
  expandedKey_5(161) <= out0_83 WHEN out0_81 = to_unsigned(16#A2#, 8) ELSE
      expandedKey_2(161);
  
  expandedKey_5(162) <= out0_83 WHEN out0_81 = to_unsigned(16#A3#, 8) ELSE
      expandedKey_2(162);
  
  expandedKey_5(163) <= out0_83 WHEN out0_81 = to_unsigned(16#A4#, 8) ELSE
      expandedKey_2(163);
  
  expandedKey_5(164) <= out0_83 WHEN out0_81 = to_unsigned(16#A5#, 8) ELSE
      expandedKey_2(164);
  
  expandedKey_5(165) <= out0_83 WHEN out0_81 = to_unsigned(16#A6#, 8) ELSE
      expandedKey_2(165);
  
  expandedKey_5(166) <= out0_83 WHEN out0_81 = to_unsigned(16#A7#, 8) ELSE
      expandedKey_2(166);
  
  expandedKey_5(167) <= out0_83 WHEN out0_81 = to_unsigned(16#A8#, 8) ELSE
      expandedKey_2(167);
  
  expandedKey_5(168) <= out0_83 WHEN out0_81 = to_unsigned(16#A9#, 8) ELSE
      expandedKey_2(168);
  
  expandedKey_5(169) <= out0_83 WHEN out0_81 = to_unsigned(16#AA#, 8) ELSE
      expandedKey_2(169);
  
  expandedKey_5(170) <= out0_83 WHEN out0_81 = to_unsigned(16#AB#, 8) ELSE
      expandedKey_2(170);
  
  expandedKey_5(171) <= out0_83 WHEN out0_81 = to_unsigned(16#AC#, 8) ELSE
      expandedKey_2(171);
  
  expandedKey_5(172) <= out0_83 WHEN out0_81 = to_unsigned(16#AD#, 8) ELSE
      expandedKey_2(172);
  
  expandedKey_5(173) <= out0_83 WHEN out0_81 = to_unsigned(16#AE#, 8) ELSE
      expandedKey_2(173);
  
  expandedKey_5(174) <= out0_83 WHEN out0_81 = to_unsigned(16#AF#, 8) ELSE
      expandedKey_2(174);
  
  expandedKey_5(175) <= out0_83 WHEN out0_81 = to_unsigned(16#B0#, 8) ELSE
      expandedKey_2(175);
  
  expandedKey_5(176) <= out0_83 WHEN out0_81 = to_unsigned(16#B1#, 8) ELSE
      expandedKey_2(176);
  
  expandedKey_5(177) <= out0_83 WHEN out0_81 = to_unsigned(16#B2#, 8) ELSE
      expandedKey_2(177);
  
  expandedKey_5(178) <= out0_83 WHEN out0_81 = to_unsigned(16#B3#, 8) ELSE
      expandedKey_2(178);
  
  expandedKey_5(179) <= out0_83 WHEN out0_81 = to_unsigned(16#B4#, 8) ELSE
      expandedKey_2(179);
  
  expandedKey_5(180) <= out0_83 WHEN out0_81 = to_unsigned(16#B5#, 8) ELSE
      expandedKey_2(180);
  
  expandedKey_5(181) <= out0_83 WHEN out0_81 = to_unsigned(16#B6#, 8) ELSE
      expandedKey_2(181);
  
  expandedKey_5(182) <= out0_83 WHEN out0_81 = to_unsigned(16#B7#, 8) ELSE
      expandedKey_2(182);
  
  expandedKey_5(183) <= out0_83 WHEN out0_81 = to_unsigned(16#B8#, 8) ELSE
      expandedKey_2(183);
  
  expandedKey_5(184) <= out0_83 WHEN out0_81 = to_unsigned(16#B9#, 8) ELSE
      expandedKey_2(184);
  
  expandedKey_5(185) <= out0_83 WHEN out0_81 = to_unsigned(16#BA#, 8) ELSE
      expandedKey_2(185);
  
  expandedKey_5(186) <= out0_83 WHEN out0_81 = to_unsigned(16#BB#, 8) ELSE
      expandedKey_2(186);
  
  expandedKey_5(187) <= out0_83 WHEN out0_81 = to_unsigned(16#BC#, 8) ELSE
      expandedKey_2(187);
  
  expandedKey_5(188) <= out0_83 WHEN out0_81 = to_unsigned(16#BD#, 8) ELSE
      expandedKey_2(188);
  
  expandedKey_5(189) <= out0_83 WHEN out0_81 = to_unsigned(16#BE#, 8) ELSE
      expandedKey_2(189);
  
  expandedKey_5(190) <= out0_83 WHEN out0_81 = to_unsigned(16#BF#, 8) ELSE
      expandedKey_2(190);
  
  expandedKey_5(191) <= out0_83 WHEN out0_81 = to_unsigned(16#C0#, 8) ELSE
      expandedKey_2(191);
  
  expandedKey_5(192) <= out0_83 WHEN out0_81 = to_unsigned(16#C1#, 8) ELSE
      expandedKey_2(192);
  
  expandedKey_5(193) <= out0_83 WHEN out0_81 = to_unsigned(16#C2#, 8) ELSE
      expandedKey_2(193);
  
  expandedKey_5(194) <= out0_83 WHEN out0_81 = to_unsigned(16#C3#, 8) ELSE
      expandedKey_2(194);
  
  expandedKey_5(195) <= out0_83 WHEN out0_81 = to_unsigned(16#C4#, 8) ELSE
      expandedKey_2(195);
  
  expandedKey_5(196) <= out0_83 WHEN out0_81 = to_unsigned(16#C5#, 8) ELSE
      expandedKey_2(196);
  
  expandedKey_5(197) <= out0_83 WHEN out0_81 = to_unsigned(16#C6#, 8) ELSE
      expandedKey_2(197);
  
  expandedKey_5(198) <= out0_83 WHEN out0_81 = to_unsigned(16#C7#, 8) ELSE
      expandedKey_2(198);
  
  expandedKey_5(199) <= out0_83 WHEN out0_81 = to_unsigned(16#C8#, 8) ELSE
      expandedKey_2(199);
  
  expandedKey_5(200) <= out0_83 WHEN out0_81 = to_unsigned(16#C9#, 8) ELSE
      expandedKey_2(200);
  
  expandedKey_5(201) <= out0_83 WHEN out0_81 = to_unsigned(16#CA#, 8) ELSE
      expandedKey_2(201);
  
  expandedKey_5(202) <= out0_83 WHEN out0_81 = to_unsigned(16#CB#, 8) ELSE
      expandedKey_2(202);
  
  expandedKey_5(203) <= out0_83 WHEN out0_81 = to_unsigned(16#CC#, 8) ELSE
      expandedKey_2(203);
  
  expandedKey_5(204) <= out0_83 WHEN out0_81 = to_unsigned(16#CD#, 8) ELSE
      expandedKey_2(204);
  
  expandedKey_5(205) <= out0_83 WHEN out0_81 = to_unsigned(16#CE#, 8) ELSE
      expandedKey_2(205);
  
  expandedKey_5(206) <= out0_83 WHEN out0_81 = to_unsigned(16#CF#, 8) ELSE
      expandedKey_2(206);
  
  expandedKey_5(207) <= out0_83 WHEN out0_81 = to_unsigned(16#D0#, 8) ELSE
      expandedKey_2(207);
  
  expandedKey_5(208) <= out0_83 WHEN out0_81 = to_unsigned(16#D1#, 8) ELSE
      expandedKey_2(208);
  
  expandedKey_5(209) <= out0_83 WHEN out0_81 = to_unsigned(16#D2#, 8) ELSE
      expandedKey_2(209);
  
  expandedKey_5(210) <= out0_83 WHEN out0_81 = to_unsigned(16#D3#, 8) ELSE
      expandedKey_2(210);
  
  expandedKey_5(211) <= out0_83 WHEN out0_81 = to_unsigned(16#D4#, 8) ELSE
      expandedKey_2(211);
  
  expandedKey_5(212) <= out0_83 WHEN out0_81 = to_unsigned(16#D5#, 8) ELSE
      expandedKey_2(212);
  
  expandedKey_5(213) <= out0_83 WHEN out0_81 = to_unsigned(16#D6#, 8) ELSE
      expandedKey_2(213);
  
  expandedKey_5(214) <= out0_83 WHEN out0_81 = to_unsigned(16#D7#, 8) ELSE
      expandedKey_2(214);
  
  expandedKey_5(215) <= out0_83 WHEN out0_81 = to_unsigned(16#D8#, 8) ELSE
      expandedKey_2(215);
  
  expandedKey_5(216) <= out0_83 WHEN out0_81 = to_unsigned(16#D9#, 8) ELSE
      expandedKey_2(216);
  
  expandedKey_5(217) <= out0_83 WHEN out0_81 = to_unsigned(16#DA#, 8) ELSE
      expandedKey_2(217);
  
  expandedKey_5(218) <= out0_83 WHEN out0_81 = to_unsigned(16#DB#, 8) ELSE
      expandedKey_2(218);
  
  expandedKey_5(219) <= out0_83 WHEN out0_81 = to_unsigned(16#DC#, 8) ELSE
      expandedKey_2(219);
  
  expandedKey_5(220) <= out0_83 WHEN out0_81 = to_unsigned(16#DD#, 8) ELSE
      expandedKey_2(220);
  
  expandedKey_5(221) <= out0_83 WHEN out0_81 = to_unsigned(16#DE#, 8) ELSE
      expandedKey_2(221);
  
  expandedKey_5(222) <= out0_83 WHEN out0_81 = to_unsigned(16#DF#, 8) ELSE
      expandedKey_2(222);
  
  expandedKey_5(223) <= out0_83 WHEN out0_81 = to_unsigned(16#E0#, 8) ELSE
      expandedKey_2(223);
  
  expandedKey_5(224) <= out0_83 WHEN out0_81 = to_unsigned(16#E1#, 8) ELSE
      expandedKey_2(224);
  
  expandedKey_5(225) <= out0_83 WHEN out0_81 = to_unsigned(16#E2#, 8) ELSE
      expandedKey_2(225);
  
  expandedKey_5(226) <= out0_83 WHEN out0_81 = to_unsigned(16#E3#, 8) ELSE
      expandedKey_2(226);
  
  expandedKey_5(227) <= out0_83 WHEN out0_81 = to_unsigned(16#E4#, 8) ELSE
      expandedKey_2(227);
  
  expandedKey_5(228) <= out0_83 WHEN out0_81 = to_unsigned(16#E5#, 8) ELSE
      expandedKey_2(228);
  
  expandedKey_5(229) <= out0_83 WHEN out0_81 = to_unsigned(16#E6#, 8) ELSE
      expandedKey_2(229);
  
  expandedKey_5(230) <= out0_83 WHEN out0_81 = to_unsigned(16#E7#, 8) ELSE
      expandedKey_2(230);
  
  expandedKey_5(231) <= out0_83 WHEN out0_81 = to_unsigned(16#E8#, 8) ELSE
      expandedKey_2(231);
  
  expandedKey_5(232) <= out0_83 WHEN out0_81 = to_unsigned(16#E9#, 8) ELSE
      expandedKey_2(232);
  
  expandedKey_5(233) <= out0_83 WHEN out0_81 = to_unsigned(16#EA#, 8) ELSE
      expandedKey_2(233);
  
  expandedKey_5(234) <= out0_83 WHEN out0_81 = to_unsigned(16#EB#, 8) ELSE
      expandedKey_2(234);
  
  expandedKey_5(235) <= out0_83 WHEN out0_81 = to_unsigned(16#EC#, 8) ELSE
      expandedKey_2(235);
  
  expandedKey_5(236) <= out0_83 WHEN out0_81 = to_unsigned(16#ED#, 8) ELSE
      expandedKey_2(236);
  
  expandedKey_5(237) <= out0_83 WHEN out0_81 = to_unsigned(16#EE#, 8) ELSE
      expandedKey_2(237);
  
  expandedKey_5(238) <= out0_83 WHEN out0_81 = to_unsigned(16#EF#, 8) ELSE
      expandedKey_2(238);
  
  expandedKey_5(239) <= out0_83 WHEN out0_81 = to_unsigned(16#F0#, 8) ELSE
      expandedKey_2(239);

  
  out0_106(0) <= expandedKey(0) WHEN out0_10 = '0' ELSE
      expandedKey(0);
  
  out0_106(1) <= expandedKey(1) WHEN out0_10 = '0' ELSE
      expandedKey(1);
  
  out0_106(2) <= expandedKey(2) WHEN out0_10 = '0' ELSE
      expandedKey(2);
  
  out0_106(3) <= expandedKey(3) WHEN out0_10 = '0' ELSE
      expandedKey(3);
  
  out0_106(4) <= expandedKey(4) WHEN out0_10 = '0' ELSE
      expandedKey(4);
  
  out0_106(5) <= expandedKey(5) WHEN out0_10 = '0' ELSE
      expandedKey(5);
  
  out0_106(6) <= expandedKey(6) WHEN out0_10 = '0' ELSE
      expandedKey(6);
  
  out0_106(7) <= expandedKey(7) WHEN out0_10 = '0' ELSE
      expandedKey(7);
  
  out0_106(8) <= expandedKey(8) WHEN out0_10 = '0' ELSE
      expandedKey(8);
  
  out0_106(9) <= expandedKey(9) WHEN out0_10 = '0' ELSE
      expandedKey(9);
  
  out0_106(10) <= expandedKey(10) WHEN out0_10 = '0' ELSE
      expandedKey(10);
  
  out0_106(11) <= expandedKey(11) WHEN out0_10 = '0' ELSE
      expandedKey(11);
  
  out0_106(12) <= expandedKey(12) WHEN out0_10 = '0' ELSE
      expandedKey(12);
  
  out0_106(13) <= expandedKey(13) WHEN out0_10 = '0' ELSE
      expandedKey(13);
  
  out0_106(14) <= expandedKey(14) WHEN out0_10 = '0' ELSE
      expandedKey(14);
  
  out0_106(15) <= expandedKey(15) WHEN out0_10 = '0' ELSE
      expandedKey(15);
  
  out0_106(16) <= expandedKey(16) WHEN out0_10 = '0' ELSE
      expandedKey(16);
  
  out0_106(17) <= expandedKey(17) WHEN out0_10 = '0' ELSE
      expandedKey(17);
  
  out0_106(18) <= expandedKey(18) WHEN out0_10 = '0' ELSE
      expandedKey(18);
  
  out0_106(19) <= expandedKey(19) WHEN out0_10 = '0' ELSE
      expandedKey(19);
  
  out0_106(20) <= expandedKey(20) WHEN out0_10 = '0' ELSE
      expandedKey(20);
  
  out0_106(21) <= expandedKey(21) WHEN out0_10 = '0' ELSE
      expandedKey(21);
  
  out0_106(22) <= expandedKey(22) WHEN out0_10 = '0' ELSE
      expandedKey(22);
  
  out0_106(23) <= expandedKey(23) WHEN out0_10 = '0' ELSE
      expandedKey(23);
  
  out0_106(24) <= expandedKey(24) WHEN out0_10 = '0' ELSE
      expandedKey(24);
  
  out0_106(25) <= expandedKey(25) WHEN out0_10 = '0' ELSE
      expandedKey(25);
  
  out0_106(26) <= expandedKey(26) WHEN out0_10 = '0' ELSE
      expandedKey(26);
  
  out0_106(27) <= expandedKey(27) WHEN out0_10 = '0' ELSE
      expandedKey(27);
  
  out0_106(28) <= expandedKey(28) WHEN out0_10 = '0' ELSE
      expandedKey(28);
  
  out0_106(29) <= expandedKey(29) WHEN out0_10 = '0' ELSE
      expandedKey(29);
  
  out0_106(30) <= expandedKey(30) WHEN out0_10 = '0' ELSE
      expandedKey(30);
  
  out0_106(31) <= expandedKey(31) WHEN out0_10 = '0' ELSE
      expandedKey(31);
  
  out0_106(32) <= expandedKey(32) WHEN out0_10 = '0' ELSE
      expandedKey(32);
  
  out0_106(33) <= expandedKey(33) WHEN out0_10 = '0' ELSE
      expandedKey(33);
  
  out0_106(34) <= expandedKey(34) WHEN out0_10 = '0' ELSE
      expandedKey(34);
  
  out0_106(35) <= expandedKey(35) WHEN out0_10 = '0' ELSE
      expandedKey(35);
  
  out0_106(36) <= expandedKey(36) WHEN out0_10 = '0' ELSE
      expandedKey(36);
  
  out0_106(37) <= expandedKey(37) WHEN out0_10 = '0' ELSE
      expandedKey(37);
  
  out0_106(38) <= expandedKey(38) WHEN out0_10 = '0' ELSE
      expandedKey(38);
  
  out0_106(39) <= expandedKey(39) WHEN out0_10 = '0' ELSE
      expandedKey(39);
  
  out0_106(40) <= expandedKey(40) WHEN out0_10 = '0' ELSE
      expandedKey(40);
  
  out0_106(41) <= expandedKey(41) WHEN out0_10 = '0' ELSE
      expandedKey(41);
  
  out0_106(42) <= expandedKey(42) WHEN out0_10 = '0' ELSE
      expandedKey(42);
  
  out0_106(43) <= expandedKey(43) WHEN out0_10 = '0' ELSE
      expandedKey(43);
  
  out0_106(44) <= expandedKey(44) WHEN out0_10 = '0' ELSE
      expandedKey(44);
  
  out0_106(45) <= expandedKey(45) WHEN out0_10 = '0' ELSE
      expandedKey(45);
  
  out0_106(46) <= expandedKey(46) WHEN out0_10 = '0' ELSE
      expandedKey(46);
  
  out0_106(47) <= expandedKey(47) WHEN out0_10 = '0' ELSE
      expandedKey(47);
  
  out0_106(48) <= expandedKey(48) WHEN out0_10 = '0' ELSE
      expandedKey(48);
  
  out0_106(49) <= expandedKey(49) WHEN out0_10 = '0' ELSE
      expandedKey(49);
  
  out0_106(50) <= expandedKey(50) WHEN out0_10 = '0' ELSE
      expandedKey(50);
  
  out0_106(51) <= expandedKey(51) WHEN out0_10 = '0' ELSE
      expandedKey(51);
  
  out0_106(52) <= expandedKey(52) WHEN out0_10 = '0' ELSE
      expandedKey(52);
  
  out0_106(53) <= expandedKey(53) WHEN out0_10 = '0' ELSE
      expandedKey(53);
  
  out0_106(54) <= expandedKey(54) WHEN out0_10 = '0' ELSE
      expandedKey(54);
  
  out0_106(55) <= expandedKey(55) WHEN out0_10 = '0' ELSE
      expandedKey(55);
  
  out0_106(56) <= expandedKey(56) WHEN out0_10 = '0' ELSE
      expandedKey(56);
  
  out0_106(57) <= expandedKey(57) WHEN out0_10 = '0' ELSE
      expandedKey(57);
  
  out0_106(58) <= expandedKey(58) WHEN out0_10 = '0' ELSE
      expandedKey(58);
  
  out0_106(59) <= expandedKey(59) WHEN out0_10 = '0' ELSE
      expandedKey(59);
  
  out0_106(60) <= expandedKey(60) WHEN out0_10 = '0' ELSE
      expandedKey(60);
  
  out0_106(61) <= expandedKey(61) WHEN out0_10 = '0' ELSE
      expandedKey(61);
  
  out0_106(62) <= expandedKey(62) WHEN out0_10 = '0' ELSE
      expandedKey(62);
  
  out0_106(63) <= expandedKey(63) WHEN out0_10 = '0' ELSE
      expandedKey(63);
  
  out0_106(64) <= expandedKey(64) WHEN out0_10 = '0' ELSE
      expandedKey(64);
  
  out0_106(65) <= expandedKey(65) WHEN out0_10 = '0' ELSE
      expandedKey(65);
  
  out0_106(66) <= expandedKey(66) WHEN out0_10 = '0' ELSE
      expandedKey(66);
  
  out0_106(67) <= expandedKey(67) WHEN out0_10 = '0' ELSE
      expandedKey(67);
  
  out0_106(68) <= expandedKey(68) WHEN out0_10 = '0' ELSE
      expandedKey(68);
  
  out0_106(69) <= expandedKey(69) WHEN out0_10 = '0' ELSE
      expandedKey(69);
  
  out0_106(70) <= expandedKey(70) WHEN out0_10 = '0' ELSE
      expandedKey(70);
  
  out0_106(71) <= expandedKey(71) WHEN out0_10 = '0' ELSE
      expandedKey(71);
  
  out0_106(72) <= expandedKey(72) WHEN out0_10 = '0' ELSE
      expandedKey(72);
  
  out0_106(73) <= expandedKey(73) WHEN out0_10 = '0' ELSE
      expandedKey(73);
  
  out0_106(74) <= expandedKey(74) WHEN out0_10 = '0' ELSE
      expandedKey(74);
  
  out0_106(75) <= expandedKey(75) WHEN out0_10 = '0' ELSE
      expandedKey(75);
  
  out0_106(76) <= expandedKey(76) WHEN out0_10 = '0' ELSE
      expandedKey(76);
  
  out0_106(77) <= expandedKey(77) WHEN out0_10 = '0' ELSE
      expandedKey(77);
  
  out0_106(78) <= expandedKey(78) WHEN out0_10 = '0' ELSE
      expandedKey(78);
  
  out0_106(79) <= expandedKey(79) WHEN out0_10 = '0' ELSE
      expandedKey(79);
  
  out0_106(80) <= expandedKey(80) WHEN out0_10 = '0' ELSE
      expandedKey(80);
  
  out0_106(81) <= expandedKey(81) WHEN out0_10 = '0' ELSE
      expandedKey(81);
  
  out0_106(82) <= expandedKey(82) WHEN out0_10 = '0' ELSE
      expandedKey(82);
  
  out0_106(83) <= expandedKey(83) WHEN out0_10 = '0' ELSE
      expandedKey(83);
  
  out0_106(84) <= expandedKey(84) WHEN out0_10 = '0' ELSE
      expandedKey(84);
  
  out0_106(85) <= expandedKey(85) WHEN out0_10 = '0' ELSE
      expandedKey(85);
  
  out0_106(86) <= expandedKey(86) WHEN out0_10 = '0' ELSE
      expandedKey(86);
  
  out0_106(87) <= expandedKey(87) WHEN out0_10 = '0' ELSE
      expandedKey(87);
  
  out0_106(88) <= expandedKey(88) WHEN out0_10 = '0' ELSE
      expandedKey(88);
  
  out0_106(89) <= expandedKey(89) WHEN out0_10 = '0' ELSE
      expandedKey(89);
  
  out0_106(90) <= expandedKey(90) WHEN out0_10 = '0' ELSE
      expandedKey(90);
  
  out0_106(91) <= expandedKey(91) WHEN out0_10 = '0' ELSE
      expandedKey(91);
  
  out0_106(92) <= expandedKey(92) WHEN out0_10 = '0' ELSE
      expandedKey(92);
  
  out0_106(93) <= expandedKey(93) WHEN out0_10 = '0' ELSE
      expandedKey(93);
  
  out0_106(94) <= expandedKey(94) WHEN out0_10 = '0' ELSE
      expandedKey(94);
  
  out0_106(95) <= expandedKey(95) WHEN out0_10 = '0' ELSE
      expandedKey(95);
  
  out0_106(96) <= expandedKey(96) WHEN out0_10 = '0' ELSE
      expandedKey(96);
  
  out0_106(97) <= expandedKey(97) WHEN out0_10 = '0' ELSE
      expandedKey(97);
  
  out0_106(98) <= expandedKey(98) WHEN out0_10 = '0' ELSE
      expandedKey(98);
  
  out0_106(99) <= expandedKey(99) WHEN out0_10 = '0' ELSE
      expandedKey(99);
  
  out0_106(100) <= expandedKey(100) WHEN out0_10 = '0' ELSE
      expandedKey(100);
  
  out0_106(101) <= expandedKey(101) WHEN out0_10 = '0' ELSE
      expandedKey(101);
  
  out0_106(102) <= expandedKey(102) WHEN out0_10 = '0' ELSE
      expandedKey(102);
  
  out0_106(103) <= expandedKey(103) WHEN out0_10 = '0' ELSE
      expandedKey(103);
  
  out0_106(104) <= expandedKey(104) WHEN out0_10 = '0' ELSE
      expandedKey(104);
  
  out0_106(105) <= expandedKey(105) WHEN out0_10 = '0' ELSE
      expandedKey(105);
  
  out0_106(106) <= expandedKey(106) WHEN out0_10 = '0' ELSE
      expandedKey(106);
  
  out0_106(107) <= expandedKey(107) WHEN out0_10 = '0' ELSE
      expandedKey(107);
  
  out0_106(108) <= expandedKey(108) WHEN out0_10 = '0' ELSE
      expandedKey(108);
  
  out0_106(109) <= expandedKey(109) WHEN out0_10 = '0' ELSE
      expandedKey(109);
  
  out0_106(110) <= expandedKey(110) WHEN out0_10 = '0' ELSE
      expandedKey(110);
  
  out0_106(111) <= expandedKey(111) WHEN out0_10 = '0' ELSE
      expandedKey(111);
  
  out0_106(112) <= expandedKey(112) WHEN out0_10 = '0' ELSE
      expandedKey(112);
  
  out0_106(113) <= expandedKey(113) WHEN out0_10 = '0' ELSE
      expandedKey(113);
  
  out0_106(114) <= expandedKey(114) WHEN out0_10 = '0' ELSE
      expandedKey(114);
  
  out0_106(115) <= expandedKey(115) WHEN out0_10 = '0' ELSE
      expandedKey(115);
  
  out0_106(116) <= expandedKey(116) WHEN out0_10 = '0' ELSE
      expandedKey(116);
  
  out0_106(117) <= expandedKey(117) WHEN out0_10 = '0' ELSE
      expandedKey(117);
  
  out0_106(118) <= expandedKey(118) WHEN out0_10 = '0' ELSE
      expandedKey(118);
  
  out0_106(119) <= expandedKey(119) WHEN out0_10 = '0' ELSE
      expandedKey(119);
  
  out0_106(120) <= expandedKey(120) WHEN out0_10 = '0' ELSE
      expandedKey(120);
  
  out0_106(121) <= expandedKey(121) WHEN out0_10 = '0' ELSE
      expandedKey(121);
  
  out0_106(122) <= expandedKey(122) WHEN out0_10 = '0' ELSE
      expandedKey(122);
  
  out0_106(123) <= expandedKey(123) WHEN out0_10 = '0' ELSE
      expandedKey(123);
  
  out0_106(124) <= expandedKey(124) WHEN out0_10 = '0' ELSE
      expandedKey(124);
  
  out0_106(125) <= expandedKey(125) WHEN out0_10 = '0' ELSE
      expandedKey(125);
  
  out0_106(126) <= expandedKey(126) WHEN out0_10 = '0' ELSE
      expandedKey(126);
  
  out0_106(127) <= expandedKey(127) WHEN out0_10 = '0' ELSE
      expandedKey(127);
  
  out0_106(128) <= expandedKey(128) WHEN out0_10 = '0' ELSE
      expandedKey(128);
  
  out0_106(129) <= expandedKey(129) WHEN out0_10 = '0' ELSE
      expandedKey(129);
  
  out0_106(130) <= expandedKey(130) WHEN out0_10 = '0' ELSE
      expandedKey(130);
  
  out0_106(131) <= expandedKey(131) WHEN out0_10 = '0' ELSE
      expandedKey(131);
  
  out0_106(132) <= expandedKey(132) WHEN out0_10 = '0' ELSE
      expandedKey(132);
  
  out0_106(133) <= expandedKey(133) WHEN out0_10 = '0' ELSE
      expandedKey(133);
  
  out0_106(134) <= expandedKey(134) WHEN out0_10 = '0' ELSE
      expandedKey(134);
  
  out0_106(135) <= expandedKey(135) WHEN out0_10 = '0' ELSE
      expandedKey(135);
  
  out0_106(136) <= expandedKey(136) WHEN out0_10 = '0' ELSE
      expandedKey(136);
  
  out0_106(137) <= expandedKey(137) WHEN out0_10 = '0' ELSE
      expandedKey(137);
  
  out0_106(138) <= expandedKey(138) WHEN out0_10 = '0' ELSE
      expandedKey(138);
  
  out0_106(139) <= expandedKey(139) WHEN out0_10 = '0' ELSE
      expandedKey(139);
  
  out0_106(140) <= expandedKey(140) WHEN out0_10 = '0' ELSE
      expandedKey(140);
  
  out0_106(141) <= expandedKey(141) WHEN out0_10 = '0' ELSE
      expandedKey(141);
  
  out0_106(142) <= expandedKey(142) WHEN out0_10 = '0' ELSE
      expandedKey(142);
  
  out0_106(143) <= expandedKey(143) WHEN out0_10 = '0' ELSE
      expandedKey(143);
  
  out0_106(144) <= expandedKey(144) WHEN out0_10 = '0' ELSE
      expandedKey(144);
  
  out0_106(145) <= expandedKey(145) WHEN out0_10 = '0' ELSE
      expandedKey(145);
  
  out0_106(146) <= expandedKey(146) WHEN out0_10 = '0' ELSE
      expandedKey(146);
  
  out0_106(147) <= expandedKey(147) WHEN out0_10 = '0' ELSE
      expandedKey(147);
  
  out0_106(148) <= expandedKey(148) WHEN out0_10 = '0' ELSE
      expandedKey(148);
  
  out0_106(149) <= expandedKey(149) WHEN out0_10 = '0' ELSE
      expandedKey(149);
  
  out0_106(150) <= expandedKey(150) WHEN out0_10 = '0' ELSE
      expandedKey(150);
  
  out0_106(151) <= expandedKey(151) WHEN out0_10 = '0' ELSE
      expandedKey(151);
  
  out0_106(152) <= expandedKey(152) WHEN out0_10 = '0' ELSE
      expandedKey(152);
  
  out0_106(153) <= expandedKey(153) WHEN out0_10 = '0' ELSE
      expandedKey(153);
  
  out0_106(154) <= expandedKey(154) WHEN out0_10 = '0' ELSE
      expandedKey(154);
  
  out0_106(155) <= expandedKey(155) WHEN out0_10 = '0' ELSE
      expandedKey(155);
  
  out0_106(156) <= expandedKey(156) WHEN out0_10 = '0' ELSE
      expandedKey(156);
  
  out0_106(157) <= expandedKey(157) WHEN out0_10 = '0' ELSE
      expandedKey(157);
  
  out0_106(158) <= expandedKey(158) WHEN out0_10 = '0' ELSE
      expandedKey(158);
  
  out0_106(159) <= expandedKey(159) WHEN out0_10 = '0' ELSE
      expandedKey(159);
  
  out0_106(160) <= expandedKey(160) WHEN out0_10 = '0' ELSE
      expandedKey(160);
  
  out0_106(161) <= expandedKey(161) WHEN out0_10 = '0' ELSE
      expandedKey(161);
  
  out0_106(162) <= expandedKey(162) WHEN out0_10 = '0' ELSE
      expandedKey(162);
  
  out0_106(163) <= expandedKey(163) WHEN out0_10 = '0' ELSE
      expandedKey(163);
  
  out0_106(164) <= expandedKey(164) WHEN out0_10 = '0' ELSE
      expandedKey(164);
  
  out0_106(165) <= expandedKey(165) WHEN out0_10 = '0' ELSE
      expandedKey(165);
  
  out0_106(166) <= expandedKey(166) WHEN out0_10 = '0' ELSE
      expandedKey(166);
  
  out0_106(167) <= expandedKey(167) WHEN out0_10 = '0' ELSE
      expandedKey(167);
  
  out0_106(168) <= expandedKey(168) WHEN out0_10 = '0' ELSE
      expandedKey(168);
  
  out0_106(169) <= expandedKey(169) WHEN out0_10 = '0' ELSE
      expandedKey(169);
  
  out0_106(170) <= expandedKey(170) WHEN out0_10 = '0' ELSE
      expandedKey(170);
  
  out0_106(171) <= expandedKey(171) WHEN out0_10 = '0' ELSE
      expandedKey(171);
  
  out0_106(172) <= expandedKey(172) WHEN out0_10 = '0' ELSE
      expandedKey(172);
  
  out0_106(173) <= expandedKey(173) WHEN out0_10 = '0' ELSE
      expandedKey(173);
  
  out0_106(174) <= expandedKey(174) WHEN out0_10 = '0' ELSE
      expandedKey(174);
  
  out0_106(175) <= expandedKey(175) WHEN out0_10 = '0' ELSE
      expandedKey(175);
  
  out0_106(176) <= expandedKey(176) WHEN out0_10 = '0' ELSE
      expandedKey(176);
  
  out0_106(177) <= expandedKey(177) WHEN out0_10 = '0' ELSE
      expandedKey(177);
  
  out0_106(178) <= expandedKey(178) WHEN out0_10 = '0' ELSE
      expandedKey(178);
  
  out0_106(179) <= expandedKey(179) WHEN out0_10 = '0' ELSE
      expandedKey(179);
  
  out0_106(180) <= expandedKey(180) WHEN out0_10 = '0' ELSE
      expandedKey(180);
  
  out0_106(181) <= expandedKey(181) WHEN out0_10 = '0' ELSE
      expandedKey(181);
  
  out0_106(182) <= expandedKey(182) WHEN out0_10 = '0' ELSE
      expandedKey(182);
  
  out0_106(183) <= expandedKey(183) WHEN out0_10 = '0' ELSE
      expandedKey(183);
  
  out0_106(184) <= expandedKey(184) WHEN out0_10 = '0' ELSE
      expandedKey(184);
  
  out0_106(185) <= expandedKey(185) WHEN out0_10 = '0' ELSE
      expandedKey(185);
  
  out0_106(186) <= expandedKey(186) WHEN out0_10 = '0' ELSE
      expandedKey(186);
  
  out0_106(187) <= expandedKey(187) WHEN out0_10 = '0' ELSE
      expandedKey(187);
  
  out0_106(188) <= expandedKey(188) WHEN out0_10 = '0' ELSE
      expandedKey(188);
  
  out0_106(189) <= expandedKey(189) WHEN out0_10 = '0' ELSE
      expandedKey(189);
  
  out0_106(190) <= expandedKey(190) WHEN out0_10 = '0' ELSE
      expandedKey(190);
  
  out0_106(191) <= expandedKey(191) WHEN out0_10 = '0' ELSE
      expandedKey(191);
  
  out0_106(192) <= expandedKey(192) WHEN out0_10 = '0' ELSE
      expandedKey(192);
  
  out0_106(193) <= expandedKey(193) WHEN out0_10 = '0' ELSE
      expandedKey(193);
  
  out0_106(194) <= expandedKey(194) WHEN out0_10 = '0' ELSE
      expandedKey(194);
  
  out0_106(195) <= expandedKey(195) WHEN out0_10 = '0' ELSE
      expandedKey(195);
  
  out0_106(196) <= expandedKey(196) WHEN out0_10 = '0' ELSE
      expandedKey(196);
  
  out0_106(197) <= expandedKey(197) WHEN out0_10 = '0' ELSE
      expandedKey(197);
  
  out0_106(198) <= expandedKey(198) WHEN out0_10 = '0' ELSE
      expandedKey(198);
  
  out0_106(199) <= expandedKey(199) WHEN out0_10 = '0' ELSE
      expandedKey(199);
  
  out0_106(200) <= expandedKey(200) WHEN out0_10 = '0' ELSE
      expandedKey(200);
  
  out0_106(201) <= expandedKey(201) WHEN out0_10 = '0' ELSE
      expandedKey(201);
  
  out0_106(202) <= expandedKey(202) WHEN out0_10 = '0' ELSE
      expandedKey(202);
  
  out0_106(203) <= expandedKey(203) WHEN out0_10 = '0' ELSE
      expandedKey(203);
  
  out0_106(204) <= expandedKey(204) WHEN out0_10 = '0' ELSE
      expandedKey(204);
  
  out0_106(205) <= expandedKey(205) WHEN out0_10 = '0' ELSE
      expandedKey(205);
  
  out0_106(206) <= expandedKey(206) WHEN out0_10 = '0' ELSE
      expandedKey(206);
  
  out0_106(207) <= expandedKey(207) WHEN out0_10 = '0' ELSE
      expandedKey(207);
  
  out0_106(208) <= expandedKey(208) WHEN out0_10 = '0' ELSE
      expandedKey(208);
  
  out0_106(209) <= expandedKey(209) WHEN out0_10 = '0' ELSE
      expandedKey(209);
  
  out0_106(210) <= expandedKey(210) WHEN out0_10 = '0' ELSE
      expandedKey(210);
  
  out0_106(211) <= expandedKey(211) WHEN out0_10 = '0' ELSE
      expandedKey(211);
  
  out0_106(212) <= expandedKey(212) WHEN out0_10 = '0' ELSE
      expandedKey(212);
  
  out0_106(213) <= expandedKey(213) WHEN out0_10 = '0' ELSE
      expandedKey(213);
  
  out0_106(214) <= expandedKey(214) WHEN out0_10 = '0' ELSE
      expandedKey(214);
  
  out0_106(215) <= expandedKey(215) WHEN out0_10 = '0' ELSE
      expandedKey(215);
  
  out0_106(216) <= expandedKey(216) WHEN out0_10 = '0' ELSE
      expandedKey(216);
  
  out0_106(217) <= expandedKey(217) WHEN out0_10 = '0' ELSE
      expandedKey(217);
  
  out0_106(218) <= expandedKey(218) WHEN out0_10 = '0' ELSE
      expandedKey(218);
  
  out0_106(219) <= expandedKey(219) WHEN out0_10 = '0' ELSE
      expandedKey(219);
  
  out0_106(220) <= expandedKey(220) WHEN out0_10 = '0' ELSE
      expandedKey(220);
  
  out0_106(221) <= expandedKey(221) WHEN out0_10 = '0' ELSE
      expandedKey(221);
  
  out0_106(222) <= expandedKey(222) WHEN out0_10 = '0' ELSE
      expandedKey(222);
  
  out0_106(223) <= expandedKey(223) WHEN out0_10 = '0' ELSE
      expandedKey(223);
  
  out0_106(224) <= expandedKey(224) WHEN out0_10 = '0' ELSE
      expandedKey(224);
  
  out0_106(225) <= expandedKey(225) WHEN out0_10 = '0' ELSE
      expandedKey(225);
  
  out0_106(226) <= expandedKey(226) WHEN out0_10 = '0' ELSE
      expandedKey(226);
  
  out0_106(227) <= expandedKey(227) WHEN out0_10 = '0' ELSE
      expandedKey(227);
  
  out0_106(228) <= expandedKey(228) WHEN out0_10 = '0' ELSE
      expandedKey(228);
  
  out0_106(229) <= expandedKey(229) WHEN out0_10 = '0' ELSE
      expandedKey(229);
  
  out0_106(230) <= expandedKey(230) WHEN out0_10 = '0' ELSE
      expandedKey(230);
  
  out0_106(231) <= expandedKey(231) WHEN out0_10 = '0' ELSE
      expandedKey(231);
  
  out0_106(232) <= expandedKey(232) WHEN out0_10 = '0' ELSE
      expandedKey(232);
  
  out0_106(233) <= expandedKey(233) WHEN out0_10 = '0' ELSE
      expandedKey(233);
  
  out0_106(234) <= expandedKey(234) WHEN out0_10 = '0' ELSE
      expandedKey(234);
  
  out0_106(235) <= expandedKey(235) WHEN out0_10 = '0' ELSE
      expandedKey(235);
  
  out0_106(236) <= expandedKey(236) WHEN out0_10 = '0' ELSE
      expandedKey(236);
  
  out0_106(237) <= expandedKey(237) WHEN out0_10 = '0' ELSE
      expandedKey(237);
  
  out0_106(238) <= expandedKey(238) WHEN out0_10 = '0' ELSE
      expandedKey(238);
  
  out0_106(239) <= expandedKey(239) WHEN out0_10 = '0' ELSE
      expandedKey(239);

  
  out0_107(0) <= out0_106(0) WHEN out0_12 = '0' ELSE
      expandedKey(0);
  
  out0_107(1) <= out0_106(1) WHEN out0_12 = '0' ELSE
      expandedKey(1);
  
  out0_107(2) <= out0_106(2) WHEN out0_12 = '0' ELSE
      expandedKey(2);
  
  out0_107(3) <= out0_106(3) WHEN out0_12 = '0' ELSE
      expandedKey(3);
  
  out0_107(4) <= out0_106(4) WHEN out0_12 = '0' ELSE
      expandedKey(4);
  
  out0_107(5) <= out0_106(5) WHEN out0_12 = '0' ELSE
      expandedKey(5);
  
  out0_107(6) <= out0_106(6) WHEN out0_12 = '0' ELSE
      expandedKey(6);
  
  out0_107(7) <= out0_106(7) WHEN out0_12 = '0' ELSE
      expandedKey(7);
  
  out0_107(8) <= out0_106(8) WHEN out0_12 = '0' ELSE
      expandedKey(8);
  
  out0_107(9) <= out0_106(9) WHEN out0_12 = '0' ELSE
      expandedKey(9);
  
  out0_107(10) <= out0_106(10) WHEN out0_12 = '0' ELSE
      expandedKey(10);
  
  out0_107(11) <= out0_106(11) WHEN out0_12 = '0' ELSE
      expandedKey(11);
  
  out0_107(12) <= out0_106(12) WHEN out0_12 = '0' ELSE
      expandedKey(12);
  
  out0_107(13) <= out0_106(13) WHEN out0_12 = '0' ELSE
      expandedKey(13);
  
  out0_107(14) <= out0_106(14) WHEN out0_12 = '0' ELSE
      expandedKey(14);
  
  out0_107(15) <= out0_106(15) WHEN out0_12 = '0' ELSE
      expandedKey(15);
  
  out0_107(16) <= out0_106(16) WHEN out0_12 = '0' ELSE
      expandedKey(16);
  
  out0_107(17) <= out0_106(17) WHEN out0_12 = '0' ELSE
      expandedKey(17);
  
  out0_107(18) <= out0_106(18) WHEN out0_12 = '0' ELSE
      expandedKey(18);
  
  out0_107(19) <= out0_106(19) WHEN out0_12 = '0' ELSE
      expandedKey(19);
  
  out0_107(20) <= out0_106(20) WHEN out0_12 = '0' ELSE
      expandedKey(20);
  
  out0_107(21) <= out0_106(21) WHEN out0_12 = '0' ELSE
      expandedKey(21);
  
  out0_107(22) <= out0_106(22) WHEN out0_12 = '0' ELSE
      expandedKey(22);
  
  out0_107(23) <= out0_106(23) WHEN out0_12 = '0' ELSE
      expandedKey(23);
  
  out0_107(24) <= out0_106(24) WHEN out0_12 = '0' ELSE
      expandedKey(24);
  
  out0_107(25) <= out0_106(25) WHEN out0_12 = '0' ELSE
      expandedKey(25);
  
  out0_107(26) <= out0_106(26) WHEN out0_12 = '0' ELSE
      expandedKey(26);
  
  out0_107(27) <= out0_106(27) WHEN out0_12 = '0' ELSE
      expandedKey(27);
  
  out0_107(28) <= out0_106(28) WHEN out0_12 = '0' ELSE
      expandedKey(28);
  
  out0_107(29) <= out0_106(29) WHEN out0_12 = '0' ELSE
      expandedKey(29);
  
  out0_107(30) <= out0_106(30) WHEN out0_12 = '0' ELSE
      expandedKey(30);
  
  out0_107(31) <= out0_106(31) WHEN out0_12 = '0' ELSE
      expandedKey(31);
  
  out0_107(32) <= out0_106(32) WHEN out0_12 = '0' ELSE
      expandedKey(32);
  
  out0_107(33) <= out0_106(33) WHEN out0_12 = '0' ELSE
      expandedKey(33);
  
  out0_107(34) <= out0_106(34) WHEN out0_12 = '0' ELSE
      expandedKey(34);
  
  out0_107(35) <= out0_106(35) WHEN out0_12 = '0' ELSE
      expandedKey(35);
  
  out0_107(36) <= out0_106(36) WHEN out0_12 = '0' ELSE
      expandedKey(36);
  
  out0_107(37) <= out0_106(37) WHEN out0_12 = '0' ELSE
      expandedKey(37);
  
  out0_107(38) <= out0_106(38) WHEN out0_12 = '0' ELSE
      expandedKey(38);
  
  out0_107(39) <= out0_106(39) WHEN out0_12 = '0' ELSE
      expandedKey(39);
  
  out0_107(40) <= out0_106(40) WHEN out0_12 = '0' ELSE
      expandedKey(40);
  
  out0_107(41) <= out0_106(41) WHEN out0_12 = '0' ELSE
      expandedKey(41);
  
  out0_107(42) <= out0_106(42) WHEN out0_12 = '0' ELSE
      expandedKey(42);
  
  out0_107(43) <= out0_106(43) WHEN out0_12 = '0' ELSE
      expandedKey(43);
  
  out0_107(44) <= out0_106(44) WHEN out0_12 = '0' ELSE
      expandedKey(44);
  
  out0_107(45) <= out0_106(45) WHEN out0_12 = '0' ELSE
      expandedKey(45);
  
  out0_107(46) <= out0_106(46) WHEN out0_12 = '0' ELSE
      expandedKey(46);
  
  out0_107(47) <= out0_106(47) WHEN out0_12 = '0' ELSE
      expandedKey(47);
  
  out0_107(48) <= out0_106(48) WHEN out0_12 = '0' ELSE
      expandedKey(48);
  
  out0_107(49) <= out0_106(49) WHEN out0_12 = '0' ELSE
      expandedKey(49);
  
  out0_107(50) <= out0_106(50) WHEN out0_12 = '0' ELSE
      expandedKey(50);
  
  out0_107(51) <= out0_106(51) WHEN out0_12 = '0' ELSE
      expandedKey(51);
  
  out0_107(52) <= out0_106(52) WHEN out0_12 = '0' ELSE
      expandedKey(52);
  
  out0_107(53) <= out0_106(53) WHEN out0_12 = '0' ELSE
      expandedKey(53);
  
  out0_107(54) <= out0_106(54) WHEN out0_12 = '0' ELSE
      expandedKey(54);
  
  out0_107(55) <= out0_106(55) WHEN out0_12 = '0' ELSE
      expandedKey(55);
  
  out0_107(56) <= out0_106(56) WHEN out0_12 = '0' ELSE
      expandedKey(56);
  
  out0_107(57) <= out0_106(57) WHEN out0_12 = '0' ELSE
      expandedKey(57);
  
  out0_107(58) <= out0_106(58) WHEN out0_12 = '0' ELSE
      expandedKey(58);
  
  out0_107(59) <= out0_106(59) WHEN out0_12 = '0' ELSE
      expandedKey(59);
  
  out0_107(60) <= out0_106(60) WHEN out0_12 = '0' ELSE
      expandedKey(60);
  
  out0_107(61) <= out0_106(61) WHEN out0_12 = '0' ELSE
      expandedKey(61);
  
  out0_107(62) <= out0_106(62) WHEN out0_12 = '0' ELSE
      expandedKey(62);
  
  out0_107(63) <= out0_106(63) WHEN out0_12 = '0' ELSE
      expandedKey(63);
  
  out0_107(64) <= out0_106(64) WHEN out0_12 = '0' ELSE
      expandedKey(64);
  
  out0_107(65) <= out0_106(65) WHEN out0_12 = '0' ELSE
      expandedKey(65);
  
  out0_107(66) <= out0_106(66) WHEN out0_12 = '0' ELSE
      expandedKey(66);
  
  out0_107(67) <= out0_106(67) WHEN out0_12 = '0' ELSE
      expandedKey(67);
  
  out0_107(68) <= out0_106(68) WHEN out0_12 = '0' ELSE
      expandedKey(68);
  
  out0_107(69) <= out0_106(69) WHEN out0_12 = '0' ELSE
      expandedKey(69);
  
  out0_107(70) <= out0_106(70) WHEN out0_12 = '0' ELSE
      expandedKey(70);
  
  out0_107(71) <= out0_106(71) WHEN out0_12 = '0' ELSE
      expandedKey(71);
  
  out0_107(72) <= out0_106(72) WHEN out0_12 = '0' ELSE
      expandedKey(72);
  
  out0_107(73) <= out0_106(73) WHEN out0_12 = '0' ELSE
      expandedKey(73);
  
  out0_107(74) <= out0_106(74) WHEN out0_12 = '0' ELSE
      expandedKey(74);
  
  out0_107(75) <= out0_106(75) WHEN out0_12 = '0' ELSE
      expandedKey(75);
  
  out0_107(76) <= out0_106(76) WHEN out0_12 = '0' ELSE
      expandedKey(76);
  
  out0_107(77) <= out0_106(77) WHEN out0_12 = '0' ELSE
      expandedKey(77);
  
  out0_107(78) <= out0_106(78) WHEN out0_12 = '0' ELSE
      expandedKey(78);
  
  out0_107(79) <= out0_106(79) WHEN out0_12 = '0' ELSE
      expandedKey(79);
  
  out0_107(80) <= out0_106(80) WHEN out0_12 = '0' ELSE
      expandedKey(80);
  
  out0_107(81) <= out0_106(81) WHEN out0_12 = '0' ELSE
      expandedKey(81);
  
  out0_107(82) <= out0_106(82) WHEN out0_12 = '0' ELSE
      expandedKey(82);
  
  out0_107(83) <= out0_106(83) WHEN out0_12 = '0' ELSE
      expandedKey(83);
  
  out0_107(84) <= out0_106(84) WHEN out0_12 = '0' ELSE
      expandedKey(84);
  
  out0_107(85) <= out0_106(85) WHEN out0_12 = '0' ELSE
      expandedKey(85);
  
  out0_107(86) <= out0_106(86) WHEN out0_12 = '0' ELSE
      expandedKey(86);
  
  out0_107(87) <= out0_106(87) WHEN out0_12 = '0' ELSE
      expandedKey(87);
  
  out0_107(88) <= out0_106(88) WHEN out0_12 = '0' ELSE
      expandedKey(88);
  
  out0_107(89) <= out0_106(89) WHEN out0_12 = '0' ELSE
      expandedKey(89);
  
  out0_107(90) <= out0_106(90) WHEN out0_12 = '0' ELSE
      expandedKey(90);
  
  out0_107(91) <= out0_106(91) WHEN out0_12 = '0' ELSE
      expandedKey(91);
  
  out0_107(92) <= out0_106(92) WHEN out0_12 = '0' ELSE
      expandedKey(92);
  
  out0_107(93) <= out0_106(93) WHEN out0_12 = '0' ELSE
      expandedKey(93);
  
  out0_107(94) <= out0_106(94) WHEN out0_12 = '0' ELSE
      expandedKey(94);
  
  out0_107(95) <= out0_106(95) WHEN out0_12 = '0' ELSE
      expandedKey(95);
  
  out0_107(96) <= out0_106(96) WHEN out0_12 = '0' ELSE
      expandedKey(96);
  
  out0_107(97) <= out0_106(97) WHEN out0_12 = '0' ELSE
      expandedKey(97);
  
  out0_107(98) <= out0_106(98) WHEN out0_12 = '0' ELSE
      expandedKey(98);
  
  out0_107(99) <= out0_106(99) WHEN out0_12 = '0' ELSE
      expandedKey(99);
  
  out0_107(100) <= out0_106(100) WHEN out0_12 = '0' ELSE
      expandedKey(100);
  
  out0_107(101) <= out0_106(101) WHEN out0_12 = '0' ELSE
      expandedKey(101);
  
  out0_107(102) <= out0_106(102) WHEN out0_12 = '0' ELSE
      expandedKey(102);
  
  out0_107(103) <= out0_106(103) WHEN out0_12 = '0' ELSE
      expandedKey(103);
  
  out0_107(104) <= out0_106(104) WHEN out0_12 = '0' ELSE
      expandedKey(104);
  
  out0_107(105) <= out0_106(105) WHEN out0_12 = '0' ELSE
      expandedKey(105);
  
  out0_107(106) <= out0_106(106) WHEN out0_12 = '0' ELSE
      expandedKey(106);
  
  out0_107(107) <= out0_106(107) WHEN out0_12 = '0' ELSE
      expandedKey(107);
  
  out0_107(108) <= out0_106(108) WHEN out0_12 = '0' ELSE
      expandedKey(108);
  
  out0_107(109) <= out0_106(109) WHEN out0_12 = '0' ELSE
      expandedKey(109);
  
  out0_107(110) <= out0_106(110) WHEN out0_12 = '0' ELSE
      expandedKey(110);
  
  out0_107(111) <= out0_106(111) WHEN out0_12 = '0' ELSE
      expandedKey(111);
  
  out0_107(112) <= out0_106(112) WHEN out0_12 = '0' ELSE
      expandedKey(112);
  
  out0_107(113) <= out0_106(113) WHEN out0_12 = '0' ELSE
      expandedKey(113);
  
  out0_107(114) <= out0_106(114) WHEN out0_12 = '0' ELSE
      expandedKey(114);
  
  out0_107(115) <= out0_106(115) WHEN out0_12 = '0' ELSE
      expandedKey(115);
  
  out0_107(116) <= out0_106(116) WHEN out0_12 = '0' ELSE
      expandedKey(116);
  
  out0_107(117) <= out0_106(117) WHEN out0_12 = '0' ELSE
      expandedKey(117);
  
  out0_107(118) <= out0_106(118) WHEN out0_12 = '0' ELSE
      expandedKey(118);
  
  out0_107(119) <= out0_106(119) WHEN out0_12 = '0' ELSE
      expandedKey(119);
  
  out0_107(120) <= out0_106(120) WHEN out0_12 = '0' ELSE
      expandedKey(120);
  
  out0_107(121) <= out0_106(121) WHEN out0_12 = '0' ELSE
      expandedKey(121);
  
  out0_107(122) <= out0_106(122) WHEN out0_12 = '0' ELSE
      expandedKey(122);
  
  out0_107(123) <= out0_106(123) WHEN out0_12 = '0' ELSE
      expandedKey(123);
  
  out0_107(124) <= out0_106(124) WHEN out0_12 = '0' ELSE
      expandedKey(124);
  
  out0_107(125) <= out0_106(125) WHEN out0_12 = '0' ELSE
      expandedKey(125);
  
  out0_107(126) <= out0_106(126) WHEN out0_12 = '0' ELSE
      expandedKey(126);
  
  out0_107(127) <= out0_106(127) WHEN out0_12 = '0' ELSE
      expandedKey(127);
  
  out0_107(128) <= out0_106(128) WHEN out0_12 = '0' ELSE
      expandedKey(128);
  
  out0_107(129) <= out0_106(129) WHEN out0_12 = '0' ELSE
      expandedKey(129);
  
  out0_107(130) <= out0_106(130) WHEN out0_12 = '0' ELSE
      expandedKey(130);
  
  out0_107(131) <= out0_106(131) WHEN out0_12 = '0' ELSE
      expandedKey(131);
  
  out0_107(132) <= out0_106(132) WHEN out0_12 = '0' ELSE
      expandedKey(132);
  
  out0_107(133) <= out0_106(133) WHEN out0_12 = '0' ELSE
      expandedKey(133);
  
  out0_107(134) <= out0_106(134) WHEN out0_12 = '0' ELSE
      expandedKey(134);
  
  out0_107(135) <= out0_106(135) WHEN out0_12 = '0' ELSE
      expandedKey(135);
  
  out0_107(136) <= out0_106(136) WHEN out0_12 = '0' ELSE
      expandedKey(136);
  
  out0_107(137) <= out0_106(137) WHEN out0_12 = '0' ELSE
      expandedKey(137);
  
  out0_107(138) <= out0_106(138) WHEN out0_12 = '0' ELSE
      expandedKey(138);
  
  out0_107(139) <= out0_106(139) WHEN out0_12 = '0' ELSE
      expandedKey(139);
  
  out0_107(140) <= out0_106(140) WHEN out0_12 = '0' ELSE
      expandedKey(140);
  
  out0_107(141) <= out0_106(141) WHEN out0_12 = '0' ELSE
      expandedKey(141);
  
  out0_107(142) <= out0_106(142) WHEN out0_12 = '0' ELSE
      expandedKey(142);
  
  out0_107(143) <= out0_106(143) WHEN out0_12 = '0' ELSE
      expandedKey(143);
  
  out0_107(144) <= out0_106(144) WHEN out0_12 = '0' ELSE
      expandedKey(144);
  
  out0_107(145) <= out0_106(145) WHEN out0_12 = '0' ELSE
      expandedKey(145);
  
  out0_107(146) <= out0_106(146) WHEN out0_12 = '0' ELSE
      expandedKey(146);
  
  out0_107(147) <= out0_106(147) WHEN out0_12 = '0' ELSE
      expandedKey(147);
  
  out0_107(148) <= out0_106(148) WHEN out0_12 = '0' ELSE
      expandedKey(148);
  
  out0_107(149) <= out0_106(149) WHEN out0_12 = '0' ELSE
      expandedKey(149);
  
  out0_107(150) <= out0_106(150) WHEN out0_12 = '0' ELSE
      expandedKey(150);
  
  out0_107(151) <= out0_106(151) WHEN out0_12 = '0' ELSE
      expandedKey(151);
  
  out0_107(152) <= out0_106(152) WHEN out0_12 = '0' ELSE
      expandedKey(152);
  
  out0_107(153) <= out0_106(153) WHEN out0_12 = '0' ELSE
      expandedKey(153);
  
  out0_107(154) <= out0_106(154) WHEN out0_12 = '0' ELSE
      expandedKey(154);
  
  out0_107(155) <= out0_106(155) WHEN out0_12 = '0' ELSE
      expandedKey(155);
  
  out0_107(156) <= out0_106(156) WHEN out0_12 = '0' ELSE
      expandedKey(156);
  
  out0_107(157) <= out0_106(157) WHEN out0_12 = '0' ELSE
      expandedKey(157);
  
  out0_107(158) <= out0_106(158) WHEN out0_12 = '0' ELSE
      expandedKey(158);
  
  out0_107(159) <= out0_106(159) WHEN out0_12 = '0' ELSE
      expandedKey(159);
  
  out0_107(160) <= out0_106(160) WHEN out0_12 = '0' ELSE
      expandedKey(160);
  
  out0_107(161) <= out0_106(161) WHEN out0_12 = '0' ELSE
      expandedKey(161);
  
  out0_107(162) <= out0_106(162) WHEN out0_12 = '0' ELSE
      expandedKey(162);
  
  out0_107(163) <= out0_106(163) WHEN out0_12 = '0' ELSE
      expandedKey(163);
  
  out0_107(164) <= out0_106(164) WHEN out0_12 = '0' ELSE
      expandedKey(164);
  
  out0_107(165) <= out0_106(165) WHEN out0_12 = '0' ELSE
      expandedKey(165);
  
  out0_107(166) <= out0_106(166) WHEN out0_12 = '0' ELSE
      expandedKey(166);
  
  out0_107(167) <= out0_106(167) WHEN out0_12 = '0' ELSE
      expandedKey(167);
  
  out0_107(168) <= out0_106(168) WHEN out0_12 = '0' ELSE
      expandedKey(168);
  
  out0_107(169) <= out0_106(169) WHEN out0_12 = '0' ELSE
      expandedKey(169);
  
  out0_107(170) <= out0_106(170) WHEN out0_12 = '0' ELSE
      expandedKey(170);
  
  out0_107(171) <= out0_106(171) WHEN out0_12 = '0' ELSE
      expandedKey(171);
  
  out0_107(172) <= out0_106(172) WHEN out0_12 = '0' ELSE
      expandedKey(172);
  
  out0_107(173) <= out0_106(173) WHEN out0_12 = '0' ELSE
      expandedKey(173);
  
  out0_107(174) <= out0_106(174) WHEN out0_12 = '0' ELSE
      expandedKey(174);
  
  out0_107(175) <= out0_106(175) WHEN out0_12 = '0' ELSE
      expandedKey(175);
  
  out0_107(176) <= out0_106(176) WHEN out0_12 = '0' ELSE
      expandedKey(176);
  
  out0_107(177) <= out0_106(177) WHEN out0_12 = '0' ELSE
      expandedKey(177);
  
  out0_107(178) <= out0_106(178) WHEN out0_12 = '0' ELSE
      expandedKey(178);
  
  out0_107(179) <= out0_106(179) WHEN out0_12 = '0' ELSE
      expandedKey(179);
  
  out0_107(180) <= out0_106(180) WHEN out0_12 = '0' ELSE
      expandedKey(180);
  
  out0_107(181) <= out0_106(181) WHEN out0_12 = '0' ELSE
      expandedKey(181);
  
  out0_107(182) <= out0_106(182) WHEN out0_12 = '0' ELSE
      expandedKey(182);
  
  out0_107(183) <= out0_106(183) WHEN out0_12 = '0' ELSE
      expandedKey(183);
  
  out0_107(184) <= out0_106(184) WHEN out0_12 = '0' ELSE
      expandedKey(184);
  
  out0_107(185) <= out0_106(185) WHEN out0_12 = '0' ELSE
      expandedKey(185);
  
  out0_107(186) <= out0_106(186) WHEN out0_12 = '0' ELSE
      expandedKey(186);
  
  out0_107(187) <= out0_106(187) WHEN out0_12 = '0' ELSE
      expandedKey(187);
  
  out0_107(188) <= out0_106(188) WHEN out0_12 = '0' ELSE
      expandedKey(188);
  
  out0_107(189) <= out0_106(189) WHEN out0_12 = '0' ELSE
      expandedKey(189);
  
  out0_107(190) <= out0_106(190) WHEN out0_12 = '0' ELSE
      expandedKey(190);
  
  out0_107(191) <= out0_106(191) WHEN out0_12 = '0' ELSE
      expandedKey(191);
  
  out0_107(192) <= out0_106(192) WHEN out0_12 = '0' ELSE
      expandedKey(192);
  
  out0_107(193) <= out0_106(193) WHEN out0_12 = '0' ELSE
      expandedKey(193);
  
  out0_107(194) <= out0_106(194) WHEN out0_12 = '0' ELSE
      expandedKey(194);
  
  out0_107(195) <= out0_106(195) WHEN out0_12 = '0' ELSE
      expandedKey(195);
  
  out0_107(196) <= out0_106(196) WHEN out0_12 = '0' ELSE
      expandedKey(196);
  
  out0_107(197) <= out0_106(197) WHEN out0_12 = '0' ELSE
      expandedKey(197);
  
  out0_107(198) <= out0_106(198) WHEN out0_12 = '0' ELSE
      expandedKey(198);
  
  out0_107(199) <= out0_106(199) WHEN out0_12 = '0' ELSE
      expandedKey(199);
  
  out0_107(200) <= out0_106(200) WHEN out0_12 = '0' ELSE
      expandedKey(200);
  
  out0_107(201) <= out0_106(201) WHEN out0_12 = '0' ELSE
      expandedKey(201);
  
  out0_107(202) <= out0_106(202) WHEN out0_12 = '0' ELSE
      expandedKey(202);
  
  out0_107(203) <= out0_106(203) WHEN out0_12 = '0' ELSE
      expandedKey(203);
  
  out0_107(204) <= out0_106(204) WHEN out0_12 = '0' ELSE
      expandedKey(204);
  
  out0_107(205) <= out0_106(205) WHEN out0_12 = '0' ELSE
      expandedKey(205);
  
  out0_107(206) <= out0_106(206) WHEN out0_12 = '0' ELSE
      expandedKey(206);
  
  out0_107(207) <= out0_106(207) WHEN out0_12 = '0' ELSE
      expandedKey(207);
  
  out0_107(208) <= out0_106(208) WHEN out0_12 = '0' ELSE
      expandedKey(208);
  
  out0_107(209) <= out0_106(209) WHEN out0_12 = '0' ELSE
      expandedKey(209);
  
  out0_107(210) <= out0_106(210) WHEN out0_12 = '0' ELSE
      expandedKey(210);
  
  out0_107(211) <= out0_106(211) WHEN out0_12 = '0' ELSE
      expandedKey(211);
  
  out0_107(212) <= out0_106(212) WHEN out0_12 = '0' ELSE
      expandedKey(212);
  
  out0_107(213) <= out0_106(213) WHEN out0_12 = '0' ELSE
      expandedKey(213);
  
  out0_107(214) <= out0_106(214) WHEN out0_12 = '0' ELSE
      expandedKey(214);
  
  out0_107(215) <= out0_106(215) WHEN out0_12 = '0' ELSE
      expandedKey(215);
  
  out0_107(216) <= out0_106(216) WHEN out0_12 = '0' ELSE
      expandedKey(216);
  
  out0_107(217) <= out0_106(217) WHEN out0_12 = '0' ELSE
      expandedKey(217);
  
  out0_107(218) <= out0_106(218) WHEN out0_12 = '0' ELSE
      expandedKey(218);
  
  out0_107(219) <= out0_106(219) WHEN out0_12 = '0' ELSE
      expandedKey(219);
  
  out0_107(220) <= out0_106(220) WHEN out0_12 = '0' ELSE
      expandedKey(220);
  
  out0_107(221) <= out0_106(221) WHEN out0_12 = '0' ELSE
      expandedKey(221);
  
  out0_107(222) <= out0_106(222) WHEN out0_12 = '0' ELSE
      expandedKey(222);
  
  out0_107(223) <= out0_106(223) WHEN out0_12 = '0' ELSE
      expandedKey(223);
  
  out0_107(224) <= out0_106(224) WHEN out0_12 = '0' ELSE
      expandedKey(224);
  
  out0_107(225) <= out0_106(225) WHEN out0_12 = '0' ELSE
      expandedKey(225);
  
  out0_107(226) <= out0_106(226) WHEN out0_12 = '0' ELSE
      expandedKey(226);
  
  out0_107(227) <= out0_106(227) WHEN out0_12 = '0' ELSE
      expandedKey(227);
  
  out0_107(228) <= out0_106(228) WHEN out0_12 = '0' ELSE
      expandedKey(228);
  
  out0_107(229) <= out0_106(229) WHEN out0_12 = '0' ELSE
      expandedKey(229);
  
  out0_107(230) <= out0_106(230) WHEN out0_12 = '0' ELSE
      expandedKey(230);
  
  out0_107(231) <= out0_106(231) WHEN out0_12 = '0' ELSE
      expandedKey(231);
  
  out0_107(232) <= out0_106(232) WHEN out0_12 = '0' ELSE
      expandedKey(232);
  
  out0_107(233) <= out0_106(233) WHEN out0_12 = '0' ELSE
      expandedKey(233);
  
  out0_107(234) <= out0_106(234) WHEN out0_12 = '0' ELSE
      expandedKey(234);
  
  out0_107(235) <= out0_106(235) WHEN out0_12 = '0' ELSE
      expandedKey(235);
  
  out0_107(236) <= out0_106(236) WHEN out0_12 = '0' ELSE
      expandedKey(236);
  
  out0_107(237) <= out0_106(237) WHEN out0_12 = '0' ELSE
      expandedKey(237);
  
  out0_107(238) <= out0_106(238) WHEN out0_12 = '0' ELSE
      expandedKey(238);
  
  out0_107(239) <= out0_106(239) WHEN out0_12 = '0' ELSE
      expandedKey(239);

  
  out0_108(0) <= out0_107(0) WHEN out0_14 = '0' ELSE
      expandedKey(0);
  
  out0_108(1) <= out0_107(1) WHEN out0_14 = '0' ELSE
      expandedKey(1);
  
  out0_108(2) <= out0_107(2) WHEN out0_14 = '0' ELSE
      expandedKey(2);
  
  out0_108(3) <= out0_107(3) WHEN out0_14 = '0' ELSE
      expandedKey(3);
  
  out0_108(4) <= out0_107(4) WHEN out0_14 = '0' ELSE
      expandedKey(4);
  
  out0_108(5) <= out0_107(5) WHEN out0_14 = '0' ELSE
      expandedKey(5);
  
  out0_108(6) <= out0_107(6) WHEN out0_14 = '0' ELSE
      expandedKey(6);
  
  out0_108(7) <= out0_107(7) WHEN out0_14 = '0' ELSE
      expandedKey(7);
  
  out0_108(8) <= out0_107(8) WHEN out0_14 = '0' ELSE
      expandedKey(8);
  
  out0_108(9) <= out0_107(9) WHEN out0_14 = '0' ELSE
      expandedKey(9);
  
  out0_108(10) <= out0_107(10) WHEN out0_14 = '0' ELSE
      expandedKey(10);
  
  out0_108(11) <= out0_107(11) WHEN out0_14 = '0' ELSE
      expandedKey(11);
  
  out0_108(12) <= out0_107(12) WHEN out0_14 = '0' ELSE
      expandedKey(12);
  
  out0_108(13) <= out0_107(13) WHEN out0_14 = '0' ELSE
      expandedKey(13);
  
  out0_108(14) <= out0_107(14) WHEN out0_14 = '0' ELSE
      expandedKey(14);
  
  out0_108(15) <= out0_107(15) WHEN out0_14 = '0' ELSE
      expandedKey(15);
  
  out0_108(16) <= out0_107(16) WHEN out0_14 = '0' ELSE
      expandedKey(16);
  
  out0_108(17) <= out0_107(17) WHEN out0_14 = '0' ELSE
      expandedKey(17);
  
  out0_108(18) <= out0_107(18) WHEN out0_14 = '0' ELSE
      expandedKey(18);
  
  out0_108(19) <= out0_107(19) WHEN out0_14 = '0' ELSE
      expandedKey(19);
  
  out0_108(20) <= out0_107(20) WHEN out0_14 = '0' ELSE
      expandedKey(20);
  
  out0_108(21) <= out0_107(21) WHEN out0_14 = '0' ELSE
      expandedKey(21);
  
  out0_108(22) <= out0_107(22) WHEN out0_14 = '0' ELSE
      expandedKey(22);
  
  out0_108(23) <= out0_107(23) WHEN out0_14 = '0' ELSE
      expandedKey(23);
  
  out0_108(24) <= out0_107(24) WHEN out0_14 = '0' ELSE
      expandedKey(24);
  
  out0_108(25) <= out0_107(25) WHEN out0_14 = '0' ELSE
      expandedKey(25);
  
  out0_108(26) <= out0_107(26) WHEN out0_14 = '0' ELSE
      expandedKey(26);
  
  out0_108(27) <= out0_107(27) WHEN out0_14 = '0' ELSE
      expandedKey(27);
  
  out0_108(28) <= out0_107(28) WHEN out0_14 = '0' ELSE
      expandedKey(28);
  
  out0_108(29) <= out0_107(29) WHEN out0_14 = '0' ELSE
      expandedKey(29);
  
  out0_108(30) <= out0_107(30) WHEN out0_14 = '0' ELSE
      expandedKey(30);
  
  out0_108(31) <= out0_107(31) WHEN out0_14 = '0' ELSE
      expandedKey(31);
  
  out0_108(32) <= out0_107(32) WHEN out0_14 = '0' ELSE
      expandedKey(32);
  
  out0_108(33) <= out0_107(33) WHEN out0_14 = '0' ELSE
      expandedKey(33);
  
  out0_108(34) <= out0_107(34) WHEN out0_14 = '0' ELSE
      expandedKey(34);
  
  out0_108(35) <= out0_107(35) WHEN out0_14 = '0' ELSE
      expandedKey(35);
  
  out0_108(36) <= out0_107(36) WHEN out0_14 = '0' ELSE
      expandedKey(36);
  
  out0_108(37) <= out0_107(37) WHEN out0_14 = '0' ELSE
      expandedKey(37);
  
  out0_108(38) <= out0_107(38) WHEN out0_14 = '0' ELSE
      expandedKey(38);
  
  out0_108(39) <= out0_107(39) WHEN out0_14 = '0' ELSE
      expandedKey(39);
  
  out0_108(40) <= out0_107(40) WHEN out0_14 = '0' ELSE
      expandedKey(40);
  
  out0_108(41) <= out0_107(41) WHEN out0_14 = '0' ELSE
      expandedKey(41);
  
  out0_108(42) <= out0_107(42) WHEN out0_14 = '0' ELSE
      expandedKey(42);
  
  out0_108(43) <= out0_107(43) WHEN out0_14 = '0' ELSE
      expandedKey(43);
  
  out0_108(44) <= out0_107(44) WHEN out0_14 = '0' ELSE
      expandedKey(44);
  
  out0_108(45) <= out0_107(45) WHEN out0_14 = '0' ELSE
      expandedKey(45);
  
  out0_108(46) <= out0_107(46) WHEN out0_14 = '0' ELSE
      expandedKey(46);
  
  out0_108(47) <= out0_107(47) WHEN out0_14 = '0' ELSE
      expandedKey(47);
  
  out0_108(48) <= out0_107(48) WHEN out0_14 = '0' ELSE
      expandedKey(48);
  
  out0_108(49) <= out0_107(49) WHEN out0_14 = '0' ELSE
      expandedKey(49);
  
  out0_108(50) <= out0_107(50) WHEN out0_14 = '0' ELSE
      expandedKey(50);
  
  out0_108(51) <= out0_107(51) WHEN out0_14 = '0' ELSE
      expandedKey(51);
  
  out0_108(52) <= out0_107(52) WHEN out0_14 = '0' ELSE
      expandedKey(52);
  
  out0_108(53) <= out0_107(53) WHEN out0_14 = '0' ELSE
      expandedKey(53);
  
  out0_108(54) <= out0_107(54) WHEN out0_14 = '0' ELSE
      expandedKey(54);
  
  out0_108(55) <= out0_107(55) WHEN out0_14 = '0' ELSE
      expandedKey(55);
  
  out0_108(56) <= out0_107(56) WHEN out0_14 = '0' ELSE
      expandedKey(56);
  
  out0_108(57) <= out0_107(57) WHEN out0_14 = '0' ELSE
      expandedKey(57);
  
  out0_108(58) <= out0_107(58) WHEN out0_14 = '0' ELSE
      expandedKey(58);
  
  out0_108(59) <= out0_107(59) WHEN out0_14 = '0' ELSE
      expandedKey(59);
  
  out0_108(60) <= out0_107(60) WHEN out0_14 = '0' ELSE
      expandedKey(60);
  
  out0_108(61) <= out0_107(61) WHEN out0_14 = '0' ELSE
      expandedKey(61);
  
  out0_108(62) <= out0_107(62) WHEN out0_14 = '0' ELSE
      expandedKey(62);
  
  out0_108(63) <= out0_107(63) WHEN out0_14 = '0' ELSE
      expandedKey(63);
  
  out0_108(64) <= out0_107(64) WHEN out0_14 = '0' ELSE
      expandedKey(64);
  
  out0_108(65) <= out0_107(65) WHEN out0_14 = '0' ELSE
      expandedKey(65);
  
  out0_108(66) <= out0_107(66) WHEN out0_14 = '0' ELSE
      expandedKey(66);
  
  out0_108(67) <= out0_107(67) WHEN out0_14 = '0' ELSE
      expandedKey(67);
  
  out0_108(68) <= out0_107(68) WHEN out0_14 = '0' ELSE
      expandedKey(68);
  
  out0_108(69) <= out0_107(69) WHEN out0_14 = '0' ELSE
      expandedKey(69);
  
  out0_108(70) <= out0_107(70) WHEN out0_14 = '0' ELSE
      expandedKey(70);
  
  out0_108(71) <= out0_107(71) WHEN out0_14 = '0' ELSE
      expandedKey(71);
  
  out0_108(72) <= out0_107(72) WHEN out0_14 = '0' ELSE
      expandedKey(72);
  
  out0_108(73) <= out0_107(73) WHEN out0_14 = '0' ELSE
      expandedKey(73);
  
  out0_108(74) <= out0_107(74) WHEN out0_14 = '0' ELSE
      expandedKey(74);
  
  out0_108(75) <= out0_107(75) WHEN out0_14 = '0' ELSE
      expandedKey(75);
  
  out0_108(76) <= out0_107(76) WHEN out0_14 = '0' ELSE
      expandedKey(76);
  
  out0_108(77) <= out0_107(77) WHEN out0_14 = '0' ELSE
      expandedKey(77);
  
  out0_108(78) <= out0_107(78) WHEN out0_14 = '0' ELSE
      expandedKey(78);
  
  out0_108(79) <= out0_107(79) WHEN out0_14 = '0' ELSE
      expandedKey(79);
  
  out0_108(80) <= out0_107(80) WHEN out0_14 = '0' ELSE
      expandedKey(80);
  
  out0_108(81) <= out0_107(81) WHEN out0_14 = '0' ELSE
      expandedKey(81);
  
  out0_108(82) <= out0_107(82) WHEN out0_14 = '0' ELSE
      expandedKey(82);
  
  out0_108(83) <= out0_107(83) WHEN out0_14 = '0' ELSE
      expandedKey(83);
  
  out0_108(84) <= out0_107(84) WHEN out0_14 = '0' ELSE
      expandedKey(84);
  
  out0_108(85) <= out0_107(85) WHEN out0_14 = '0' ELSE
      expandedKey(85);
  
  out0_108(86) <= out0_107(86) WHEN out0_14 = '0' ELSE
      expandedKey(86);
  
  out0_108(87) <= out0_107(87) WHEN out0_14 = '0' ELSE
      expandedKey(87);
  
  out0_108(88) <= out0_107(88) WHEN out0_14 = '0' ELSE
      expandedKey(88);
  
  out0_108(89) <= out0_107(89) WHEN out0_14 = '0' ELSE
      expandedKey(89);
  
  out0_108(90) <= out0_107(90) WHEN out0_14 = '0' ELSE
      expandedKey(90);
  
  out0_108(91) <= out0_107(91) WHEN out0_14 = '0' ELSE
      expandedKey(91);
  
  out0_108(92) <= out0_107(92) WHEN out0_14 = '0' ELSE
      expandedKey(92);
  
  out0_108(93) <= out0_107(93) WHEN out0_14 = '0' ELSE
      expandedKey(93);
  
  out0_108(94) <= out0_107(94) WHEN out0_14 = '0' ELSE
      expandedKey(94);
  
  out0_108(95) <= out0_107(95) WHEN out0_14 = '0' ELSE
      expandedKey(95);
  
  out0_108(96) <= out0_107(96) WHEN out0_14 = '0' ELSE
      expandedKey(96);
  
  out0_108(97) <= out0_107(97) WHEN out0_14 = '0' ELSE
      expandedKey(97);
  
  out0_108(98) <= out0_107(98) WHEN out0_14 = '0' ELSE
      expandedKey(98);
  
  out0_108(99) <= out0_107(99) WHEN out0_14 = '0' ELSE
      expandedKey(99);
  
  out0_108(100) <= out0_107(100) WHEN out0_14 = '0' ELSE
      expandedKey(100);
  
  out0_108(101) <= out0_107(101) WHEN out0_14 = '0' ELSE
      expandedKey(101);
  
  out0_108(102) <= out0_107(102) WHEN out0_14 = '0' ELSE
      expandedKey(102);
  
  out0_108(103) <= out0_107(103) WHEN out0_14 = '0' ELSE
      expandedKey(103);
  
  out0_108(104) <= out0_107(104) WHEN out0_14 = '0' ELSE
      expandedKey(104);
  
  out0_108(105) <= out0_107(105) WHEN out0_14 = '0' ELSE
      expandedKey(105);
  
  out0_108(106) <= out0_107(106) WHEN out0_14 = '0' ELSE
      expandedKey(106);
  
  out0_108(107) <= out0_107(107) WHEN out0_14 = '0' ELSE
      expandedKey(107);
  
  out0_108(108) <= out0_107(108) WHEN out0_14 = '0' ELSE
      expandedKey(108);
  
  out0_108(109) <= out0_107(109) WHEN out0_14 = '0' ELSE
      expandedKey(109);
  
  out0_108(110) <= out0_107(110) WHEN out0_14 = '0' ELSE
      expandedKey(110);
  
  out0_108(111) <= out0_107(111) WHEN out0_14 = '0' ELSE
      expandedKey(111);
  
  out0_108(112) <= out0_107(112) WHEN out0_14 = '0' ELSE
      expandedKey(112);
  
  out0_108(113) <= out0_107(113) WHEN out0_14 = '0' ELSE
      expandedKey(113);
  
  out0_108(114) <= out0_107(114) WHEN out0_14 = '0' ELSE
      expandedKey(114);
  
  out0_108(115) <= out0_107(115) WHEN out0_14 = '0' ELSE
      expandedKey(115);
  
  out0_108(116) <= out0_107(116) WHEN out0_14 = '0' ELSE
      expandedKey(116);
  
  out0_108(117) <= out0_107(117) WHEN out0_14 = '0' ELSE
      expandedKey(117);
  
  out0_108(118) <= out0_107(118) WHEN out0_14 = '0' ELSE
      expandedKey(118);
  
  out0_108(119) <= out0_107(119) WHEN out0_14 = '0' ELSE
      expandedKey(119);
  
  out0_108(120) <= out0_107(120) WHEN out0_14 = '0' ELSE
      expandedKey(120);
  
  out0_108(121) <= out0_107(121) WHEN out0_14 = '0' ELSE
      expandedKey(121);
  
  out0_108(122) <= out0_107(122) WHEN out0_14 = '0' ELSE
      expandedKey(122);
  
  out0_108(123) <= out0_107(123) WHEN out0_14 = '0' ELSE
      expandedKey(123);
  
  out0_108(124) <= out0_107(124) WHEN out0_14 = '0' ELSE
      expandedKey(124);
  
  out0_108(125) <= out0_107(125) WHEN out0_14 = '0' ELSE
      expandedKey(125);
  
  out0_108(126) <= out0_107(126) WHEN out0_14 = '0' ELSE
      expandedKey(126);
  
  out0_108(127) <= out0_107(127) WHEN out0_14 = '0' ELSE
      expandedKey(127);
  
  out0_108(128) <= out0_107(128) WHEN out0_14 = '0' ELSE
      expandedKey(128);
  
  out0_108(129) <= out0_107(129) WHEN out0_14 = '0' ELSE
      expandedKey(129);
  
  out0_108(130) <= out0_107(130) WHEN out0_14 = '0' ELSE
      expandedKey(130);
  
  out0_108(131) <= out0_107(131) WHEN out0_14 = '0' ELSE
      expandedKey(131);
  
  out0_108(132) <= out0_107(132) WHEN out0_14 = '0' ELSE
      expandedKey(132);
  
  out0_108(133) <= out0_107(133) WHEN out0_14 = '0' ELSE
      expandedKey(133);
  
  out0_108(134) <= out0_107(134) WHEN out0_14 = '0' ELSE
      expandedKey(134);
  
  out0_108(135) <= out0_107(135) WHEN out0_14 = '0' ELSE
      expandedKey(135);
  
  out0_108(136) <= out0_107(136) WHEN out0_14 = '0' ELSE
      expandedKey(136);
  
  out0_108(137) <= out0_107(137) WHEN out0_14 = '0' ELSE
      expandedKey(137);
  
  out0_108(138) <= out0_107(138) WHEN out0_14 = '0' ELSE
      expandedKey(138);
  
  out0_108(139) <= out0_107(139) WHEN out0_14 = '0' ELSE
      expandedKey(139);
  
  out0_108(140) <= out0_107(140) WHEN out0_14 = '0' ELSE
      expandedKey(140);
  
  out0_108(141) <= out0_107(141) WHEN out0_14 = '0' ELSE
      expandedKey(141);
  
  out0_108(142) <= out0_107(142) WHEN out0_14 = '0' ELSE
      expandedKey(142);
  
  out0_108(143) <= out0_107(143) WHEN out0_14 = '0' ELSE
      expandedKey(143);
  
  out0_108(144) <= out0_107(144) WHEN out0_14 = '0' ELSE
      expandedKey(144);
  
  out0_108(145) <= out0_107(145) WHEN out0_14 = '0' ELSE
      expandedKey(145);
  
  out0_108(146) <= out0_107(146) WHEN out0_14 = '0' ELSE
      expandedKey(146);
  
  out0_108(147) <= out0_107(147) WHEN out0_14 = '0' ELSE
      expandedKey(147);
  
  out0_108(148) <= out0_107(148) WHEN out0_14 = '0' ELSE
      expandedKey(148);
  
  out0_108(149) <= out0_107(149) WHEN out0_14 = '0' ELSE
      expandedKey(149);
  
  out0_108(150) <= out0_107(150) WHEN out0_14 = '0' ELSE
      expandedKey(150);
  
  out0_108(151) <= out0_107(151) WHEN out0_14 = '0' ELSE
      expandedKey(151);
  
  out0_108(152) <= out0_107(152) WHEN out0_14 = '0' ELSE
      expandedKey(152);
  
  out0_108(153) <= out0_107(153) WHEN out0_14 = '0' ELSE
      expandedKey(153);
  
  out0_108(154) <= out0_107(154) WHEN out0_14 = '0' ELSE
      expandedKey(154);
  
  out0_108(155) <= out0_107(155) WHEN out0_14 = '0' ELSE
      expandedKey(155);
  
  out0_108(156) <= out0_107(156) WHEN out0_14 = '0' ELSE
      expandedKey(156);
  
  out0_108(157) <= out0_107(157) WHEN out0_14 = '0' ELSE
      expandedKey(157);
  
  out0_108(158) <= out0_107(158) WHEN out0_14 = '0' ELSE
      expandedKey(158);
  
  out0_108(159) <= out0_107(159) WHEN out0_14 = '0' ELSE
      expandedKey(159);
  
  out0_108(160) <= out0_107(160) WHEN out0_14 = '0' ELSE
      expandedKey(160);
  
  out0_108(161) <= out0_107(161) WHEN out0_14 = '0' ELSE
      expandedKey(161);
  
  out0_108(162) <= out0_107(162) WHEN out0_14 = '0' ELSE
      expandedKey(162);
  
  out0_108(163) <= out0_107(163) WHEN out0_14 = '0' ELSE
      expandedKey(163);
  
  out0_108(164) <= out0_107(164) WHEN out0_14 = '0' ELSE
      expandedKey(164);
  
  out0_108(165) <= out0_107(165) WHEN out0_14 = '0' ELSE
      expandedKey(165);
  
  out0_108(166) <= out0_107(166) WHEN out0_14 = '0' ELSE
      expandedKey(166);
  
  out0_108(167) <= out0_107(167) WHEN out0_14 = '0' ELSE
      expandedKey(167);
  
  out0_108(168) <= out0_107(168) WHEN out0_14 = '0' ELSE
      expandedKey(168);
  
  out0_108(169) <= out0_107(169) WHEN out0_14 = '0' ELSE
      expandedKey(169);
  
  out0_108(170) <= out0_107(170) WHEN out0_14 = '0' ELSE
      expandedKey(170);
  
  out0_108(171) <= out0_107(171) WHEN out0_14 = '0' ELSE
      expandedKey(171);
  
  out0_108(172) <= out0_107(172) WHEN out0_14 = '0' ELSE
      expandedKey(172);
  
  out0_108(173) <= out0_107(173) WHEN out0_14 = '0' ELSE
      expandedKey(173);
  
  out0_108(174) <= out0_107(174) WHEN out0_14 = '0' ELSE
      expandedKey(174);
  
  out0_108(175) <= out0_107(175) WHEN out0_14 = '0' ELSE
      expandedKey(175);
  
  out0_108(176) <= out0_107(176) WHEN out0_14 = '0' ELSE
      expandedKey(176);
  
  out0_108(177) <= out0_107(177) WHEN out0_14 = '0' ELSE
      expandedKey(177);
  
  out0_108(178) <= out0_107(178) WHEN out0_14 = '0' ELSE
      expandedKey(178);
  
  out0_108(179) <= out0_107(179) WHEN out0_14 = '0' ELSE
      expandedKey(179);
  
  out0_108(180) <= out0_107(180) WHEN out0_14 = '0' ELSE
      expandedKey(180);
  
  out0_108(181) <= out0_107(181) WHEN out0_14 = '0' ELSE
      expandedKey(181);
  
  out0_108(182) <= out0_107(182) WHEN out0_14 = '0' ELSE
      expandedKey(182);
  
  out0_108(183) <= out0_107(183) WHEN out0_14 = '0' ELSE
      expandedKey(183);
  
  out0_108(184) <= out0_107(184) WHEN out0_14 = '0' ELSE
      expandedKey(184);
  
  out0_108(185) <= out0_107(185) WHEN out0_14 = '0' ELSE
      expandedKey(185);
  
  out0_108(186) <= out0_107(186) WHEN out0_14 = '0' ELSE
      expandedKey(186);
  
  out0_108(187) <= out0_107(187) WHEN out0_14 = '0' ELSE
      expandedKey(187);
  
  out0_108(188) <= out0_107(188) WHEN out0_14 = '0' ELSE
      expandedKey(188);
  
  out0_108(189) <= out0_107(189) WHEN out0_14 = '0' ELSE
      expandedKey(189);
  
  out0_108(190) <= out0_107(190) WHEN out0_14 = '0' ELSE
      expandedKey(190);
  
  out0_108(191) <= out0_107(191) WHEN out0_14 = '0' ELSE
      expandedKey(191);
  
  out0_108(192) <= out0_107(192) WHEN out0_14 = '0' ELSE
      expandedKey(192);
  
  out0_108(193) <= out0_107(193) WHEN out0_14 = '0' ELSE
      expandedKey(193);
  
  out0_108(194) <= out0_107(194) WHEN out0_14 = '0' ELSE
      expandedKey(194);
  
  out0_108(195) <= out0_107(195) WHEN out0_14 = '0' ELSE
      expandedKey(195);
  
  out0_108(196) <= out0_107(196) WHEN out0_14 = '0' ELSE
      expandedKey(196);
  
  out0_108(197) <= out0_107(197) WHEN out0_14 = '0' ELSE
      expandedKey(197);
  
  out0_108(198) <= out0_107(198) WHEN out0_14 = '0' ELSE
      expandedKey(198);
  
  out0_108(199) <= out0_107(199) WHEN out0_14 = '0' ELSE
      expandedKey(199);
  
  out0_108(200) <= out0_107(200) WHEN out0_14 = '0' ELSE
      expandedKey(200);
  
  out0_108(201) <= out0_107(201) WHEN out0_14 = '0' ELSE
      expandedKey(201);
  
  out0_108(202) <= out0_107(202) WHEN out0_14 = '0' ELSE
      expandedKey(202);
  
  out0_108(203) <= out0_107(203) WHEN out0_14 = '0' ELSE
      expandedKey(203);
  
  out0_108(204) <= out0_107(204) WHEN out0_14 = '0' ELSE
      expandedKey(204);
  
  out0_108(205) <= out0_107(205) WHEN out0_14 = '0' ELSE
      expandedKey(205);
  
  out0_108(206) <= out0_107(206) WHEN out0_14 = '0' ELSE
      expandedKey(206);
  
  out0_108(207) <= out0_107(207) WHEN out0_14 = '0' ELSE
      expandedKey(207);
  
  out0_108(208) <= out0_107(208) WHEN out0_14 = '0' ELSE
      expandedKey(208);
  
  out0_108(209) <= out0_107(209) WHEN out0_14 = '0' ELSE
      expandedKey(209);
  
  out0_108(210) <= out0_107(210) WHEN out0_14 = '0' ELSE
      expandedKey(210);
  
  out0_108(211) <= out0_107(211) WHEN out0_14 = '0' ELSE
      expandedKey(211);
  
  out0_108(212) <= out0_107(212) WHEN out0_14 = '0' ELSE
      expandedKey(212);
  
  out0_108(213) <= out0_107(213) WHEN out0_14 = '0' ELSE
      expandedKey(213);
  
  out0_108(214) <= out0_107(214) WHEN out0_14 = '0' ELSE
      expandedKey(214);
  
  out0_108(215) <= out0_107(215) WHEN out0_14 = '0' ELSE
      expandedKey(215);
  
  out0_108(216) <= out0_107(216) WHEN out0_14 = '0' ELSE
      expandedKey(216);
  
  out0_108(217) <= out0_107(217) WHEN out0_14 = '0' ELSE
      expandedKey(217);
  
  out0_108(218) <= out0_107(218) WHEN out0_14 = '0' ELSE
      expandedKey(218);
  
  out0_108(219) <= out0_107(219) WHEN out0_14 = '0' ELSE
      expandedKey(219);
  
  out0_108(220) <= out0_107(220) WHEN out0_14 = '0' ELSE
      expandedKey(220);
  
  out0_108(221) <= out0_107(221) WHEN out0_14 = '0' ELSE
      expandedKey(221);
  
  out0_108(222) <= out0_107(222) WHEN out0_14 = '0' ELSE
      expandedKey(222);
  
  out0_108(223) <= out0_107(223) WHEN out0_14 = '0' ELSE
      expandedKey(223);
  
  out0_108(224) <= out0_107(224) WHEN out0_14 = '0' ELSE
      expandedKey(224);
  
  out0_108(225) <= out0_107(225) WHEN out0_14 = '0' ELSE
      expandedKey(225);
  
  out0_108(226) <= out0_107(226) WHEN out0_14 = '0' ELSE
      expandedKey(226);
  
  out0_108(227) <= out0_107(227) WHEN out0_14 = '0' ELSE
      expandedKey(227);
  
  out0_108(228) <= out0_107(228) WHEN out0_14 = '0' ELSE
      expandedKey(228);
  
  out0_108(229) <= out0_107(229) WHEN out0_14 = '0' ELSE
      expandedKey(229);
  
  out0_108(230) <= out0_107(230) WHEN out0_14 = '0' ELSE
      expandedKey(230);
  
  out0_108(231) <= out0_107(231) WHEN out0_14 = '0' ELSE
      expandedKey(231);
  
  out0_108(232) <= out0_107(232) WHEN out0_14 = '0' ELSE
      expandedKey(232);
  
  out0_108(233) <= out0_107(233) WHEN out0_14 = '0' ELSE
      expandedKey(233);
  
  out0_108(234) <= out0_107(234) WHEN out0_14 = '0' ELSE
      expandedKey(234);
  
  out0_108(235) <= out0_107(235) WHEN out0_14 = '0' ELSE
      expandedKey(235);
  
  out0_108(236) <= out0_107(236) WHEN out0_14 = '0' ELSE
      expandedKey(236);
  
  out0_108(237) <= out0_107(237) WHEN out0_14 = '0' ELSE
      expandedKey(237);
  
  out0_108(238) <= out0_107(238) WHEN out0_14 = '0' ELSE
      expandedKey(238);
  
  out0_108(239) <= out0_107(239) WHEN out0_14 = '0' ELSE
      expandedKey(239);

  
  out0_109(0) <= out0_108(0) WHEN out0_16 = '0' ELSE
      expandedKey(0);
  
  out0_109(1) <= out0_108(1) WHEN out0_16 = '0' ELSE
      expandedKey(1);
  
  out0_109(2) <= out0_108(2) WHEN out0_16 = '0' ELSE
      expandedKey(2);
  
  out0_109(3) <= out0_108(3) WHEN out0_16 = '0' ELSE
      expandedKey(3);
  
  out0_109(4) <= out0_108(4) WHEN out0_16 = '0' ELSE
      expandedKey(4);
  
  out0_109(5) <= out0_108(5) WHEN out0_16 = '0' ELSE
      expandedKey(5);
  
  out0_109(6) <= out0_108(6) WHEN out0_16 = '0' ELSE
      expandedKey(6);
  
  out0_109(7) <= out0_108(7) WHEN out0_16 = '0' ELSE
      expandedKey(7);
  
  out0_109(8) <= out0_108(8) WHEN out0_16 = '0' ELSE
      expandedKey(8);
  
  out0_109(9) <= out0_108(9) WHEN out0_16 = '0' ELSE
      expandedKey(9);
  
  out0_109(10) <= out0_108(10) WHEN out0_16 = '0' ELSE
      expandedKey(10);
  
  out0_109(11) <= out0_108(11) WHEN out0_16 = '0' ELSE
      expandedKey(11);
  
  out0_109(12) <= out0_108(12) WHEN out0_16 = '0' ELSE
      expandedKey(12);
  
  out0_109(13) <= out0_108(13) WHEN out0_16 = '0' ELSE
      expandedKey(13);
  
  out0_109(14) <= out0_108(14) WHEN out0_16 = '0' ELSE
      expandedKey(14);
  
  out0_109(15) <= out0_108(15) WHEN out0_16 = '0' ELSE
      expandedKey(15);
  
  out0_109(16) <= out0_108(16) WHEN out0_16 = '0' ELSE
      expandedKey(16);
  
  out0_109(17) <= out0_108(17) WHEN out0_16 = '0' ELSE
      expandedKey(17);
  
  out0_109(18) <= out0_108(18) WHEN out0_16 = '0' ELSE
      expandedKey(18);
  
  out0_109(19) <= out0_108(19) WHEN out0_16 = '0' ELSE
      expandedKey(19);
  
  out0_109(20) <= out0_108(20) WHEN out0_16 = '0' ELSE
      expandedKey(20);
  
  out0_109(21) <= out0_108(21) WHEN out0_16 = '0' ELSE
      expandedKey(21);
  
  out0_109(22) <= out0_108(22) WHEN out0_16 = '0' ELSE
      expandedKey(22);
  
  out0_109(23) <= out0_108(23) WHEN out0_16 = '0' ELSE
      expandedKey(23);
  
  out0_109(24) <= out0_108(24) WHEN out0_16 = '0' ELSE
      expandedKey(24);
  
  out0_109(25) <= out0_108(25) WHEN out0_16 = '0' ELSE
      expandedKey(25);
  
  out0_109(26) <= out0_108(26) WHEN out0_16 = '0' ELSE
      expandedKey(26);
  
  out0_109(27) <= out0_108(27) WHEN out0_16 = '0' ELSE
      expandedKey(27);
  
  out0_109(28) <= out0_108(28) WHEN out0_16 = '0' ELSE
      expandedKey(28);
  
  out0_109(29) <= out0_108(29) WHEN out0_16 = '0' ELSE
      expandedKey(29);
  
  out0_109(30) <= out0_108(30) WHEN out0_16 = '0' ELSE
      expandedKey(30);
  
  out0_109(31) <= out0_108(31) WHEN out0_16 = '0' ELSE
      expandedKey(31);
  
  out0_109(32) <= out0_108(32) WHEN out0_16 = '0' ELSE
      expandedKey(32);
  
  out0_109(33) <= out0_108(33) WHEN out0_16 = '0' ELSE
      expandedKey(33);
  
  out0_109(34) <= out0_108(34) WHEN out0_16 = '0' ELSE
      expandedKey(34);
  
  out0_109(35) <= out0_108(35) WHEN out0_16 = '0' ELSE
      expandedKey(35);
  
  out0_109(36) <= out0_108(36) WHEN out0_16 = '0' ELSE
      expandedKey(36);
  
  out0_109(37) <= out0_108(37) WHEN out0_16 = '0' ELSE
      expandedKey(37);
  
  out0_109(38) <= out0_108(38) WHEN out0_16 = '0' ELSE
      expandedKey(38);
  
  out0_109(39) <= out0_108(39) WHEN out0_16 = '0' ELSE
      expandedKey(39);
  
  out0_109(40) <= out0_108(40) WHEN out0_16 = '0' ELSE
      expandedKey(40);
  
  out0_109(41) <= out0_108(41) WHEN out0_16 = '0' ELSE
      expandedKey(41);
  
  out0_109(42) <= out0_108(42) WHEN out0_16 = '0' ELSE
      expandedKey(42);
  
  out0_109(43) <= out0_108(43) WHEN out0_16 = '0' ELSE
      expandedKey(43);
  
  out0_109(44) <= out0_108(44) WHEN out0_16 = '0' ELSE
      expandedKey(44);
  
  out0_109(45) <= out0_108(45) WHEN out0_16 = '0' ELSE
      expandedKey(45);
  
  out0_109(46) <= out0_108(46) WHEN out0_16 = '0' ELSE
      expandedKey(46);
  
  out0_109(47) <= out0_108(47) WHEN out0_16 = '0' ELSE
      expandedKey(47);
  
  out0_109(48) <= out0_108(48) WHEN out0_16 = '0' ELSE
      expandedKey(48);
  
  out0_109(49) <= out0_108(49) WHEN out0_16 = '0' ELSE
      expandedKey(49);
  
  out0_109(50) <= out0_108(50) WHEN out0_16 = '0' ELSE
      expandedKey(50);
  
  out0_109(51) <= out0_108(51) WHEN out0_16 = '0' ELSE
      expandedKey(51);
  
  out0_109(52) <= out0_108(52) WHEN out0_16 = '0' ELSE
      expandedKey(52);
  
  out0_109(53) <= out0_108(53) WHEN out0_16 = '0' ELSE
      expandedKey(53);
  
  out0_109(54) <= out0_108(54) WHEN out0_16 = '0' ELSE
      expandedKey(54);
  
  out0_109(55) <= out0_108(55) WHEN out0_16 = '0' ELSE
      expandedKey(55);
  
  out0_109(56) <= out0_108(56) WHEN out0_16 = '0' ELSE
      expandedKey(56);
  
  out0_109(57) <= out0_108(57) WHEN out0_16 = '0' ELSE
      expandedKey(57);
  
  out0_109(58) <= out0_108(58) WHEN out0_16 = '0' ELSE
      expandedKey(58);
  
  out0_109(59) <= out0_108(59) WHEN out0_16 = '0' ELSE
      expandedKey(59);
  
  out0_109(60) <= out0_108(60) WHEN out0_16 = '0' ELSE
      expandedKey(60);
  
  out0_109(61) <= out0_108(61) WHEN out0_16 = '0' ELSE
      expandedKey(61);
  
  out0_109(62) <= out0_108(62) WHEN out0_16 = '0' ELSE
      expandedKey(62);
  
  out0_109(63) <= out0_108(63) WHEN out0_16 = '0' ELSE
      expandedKey(63);
  
  out0_109(64) <= out0_108(64) WHEN out0_16 = '0' ELSE
      expandedKey(64);
  
  out0_109(65) <= out0_108(65) WHEN out0_16 = '0' ELSE
      expandedKey(65);
  
  out0_109(66) <= out0_108(66) WHEN out0_16 = '0' ELSE
      expandedKey(66);
  
  out0_109(67) <= out0_108(67) WHEN out0_16 = '0' ELSE
      expandedKey(67);
  
  out0_109(68) <= out0_108(68) WHEN out0_16 = '0' ELSE
      expandedKey(68);
  
  out0_109(69) <= out0_108(69) WHEN out0_16 = '0' ELSE
      expandedKey(69);
  
  out0_109(70) <= out0_108(70) WHEN out0_16 = '0' ELSE
      expandedKey(70);
  
  out0_109(71) <= out0_108(71) WHEN out0_16 = '0' ELSE
      expandedKey(71);
  
  out0_109(72) <= out0_108(72) WHEN out0_16 = '0' ELSE
      expandedKey(72);
  
  out0_109(73) <= out0_108(73) WHEN out0_16 = '0' ELSE
      expandedKey(73);
  
  out0_109(74) <= out0_108(74) WHEN out0_16 = '0' ELSE
      expandedKey(74);
  
  out0_109(75) <= out0_108(75) WHEN out0_16 = '0' ELSE
      expandedKey(75);
  
  out0_109(76) <= out0_108(76) WHEN out0_16 = '0' ELSE
      expandedKey(76);
  
  out0_109(77) <= out0_108(77) WHEN out0_16 = '0' ELSE
      expandedKey(77);
  
  out0_109(78) <= out0_108(78) WHEN out0_16 = '0' ELSE
      expandedKey(78);
  
  out0_109(79) <= out0_108(79) WHEN out0_16 = '0' ELSE
      expandedKey(79);
  
  out0_109(80) <= out0_108(80) WHEN out0_16 = '0' ELSE
      expandedKey(80);
  
  out0_109(81) <= out0_108(81) WHEN out0_16 = '0' ELSE
      expandedKey(81);
  
  out0_109(82) <= out0_108(82) WHEN out0_16 = '0' ELSE
      expandedKey(82);
  
  out0_109(83) <= out0_108(83) WHEN out0_16 = '0' ELSE
      expandedKey(83);
  
  out0_109(84) <= out0_108(84) WHEN out0_16 = '0' ELSE
      expandedKey(84);
  
  out0_109(85) <= out0_108(85) WHEN out0_16 = '0' ELSE
      expandedKey(85);
  
  out0_109(86) <= out0_108(86) WHEN out0_16 = '0' ELSE
      expandedKey(86);
  
  out0_109(87) <= out0_108(87) WHEN out0_16 = '0' ELSE
      expandedKey(87);
  
  out0_109(88) <= out0_108(88) WHEN out0_16 = '0' ELSE
      expandedKey(88);
  
  out0_109(89) <= out0_108(89) WHEN out0_16 = '0' ELSE
      expandedKey(89);
  
  out0_109(90) <= out0_108(90) WHEN out0_16 = '0' ELSE
      expandedKey(90);
  
  out0_109(91) <= out0_108(91) WHEN out0_16 = '0' ELSE
      expandedKey(91);
  
  out0_109(92) <= out0_108(92) WHEN out0_16 = '0' ELSE
      expandedKey(92);
  
  out0_109(93) <= out0_108(93) WHEN out0_16 = '0' ELSE
      expandedKey(93);
  
  out0_109(94) <= out0_108(94) WHEN out0_16 = '0' ELSE
      expandedKey(94);
  
  out0_109(95) <= out0_108(95) WHEN out0_16 = '0' ELSE
      expandedKey(95);
  
  out0_109(96) <= out0_108(96) WHEN out0_16 = '0' ELSE
      expandedKey(96);
  
  out0_109(97) <= out0_108(97) WHEN out0_16 = '0' ELSE
      expandedKey(97);
  
  out0_109(98) <= out0_108(98) WHEN out0_16 = '0' ELSE
      expandedKey(98);
  
  out0_109(99) <= out0_108(99) WHEN out0_16 = '0' ELSE
      expandedKey(99);
  
  out0_109(100) <= out0_108(100) WHEN out0_16 = '0' ELSE
      expandedKey(100);
  
  out0_109(101) <= out0_108(101) WHEN out0_16 = '0' ELSE
      expandedKey(101);
  
  out0_109(102) <= out0_108(102) WHEN out0_16 = '0' ELSE
      expandedKey(102);
  
  out0_109(103) <= out0_108(103) WHEN out0_16 = '0' ELSE
      expandedKey(103);
  
  out0_109(104) <= out0_108(104) WHEN out0_16 = '0' ELSE
      expandedKey(104);
  
  out0_109(105) <= out0_108(105) WHEN out0_16 = '0' ELSE
      expandedKey(105);
  
  out0_109(106) <= out0_108(106) WHEN out0_16 = '0' ELSE
      expandedKey(106);
  
  out0_109(107) <= out0_108(107) WHEN out0_16 = '0' ELSE
      expandedKey(107);
  
  out0_109(108) <= out0_108(108) WHEN out0_16 = '0' ELSE
      expandedKey(108);
  
  out0_109(109) <= out0_108(109) WHEN out0_16 = '0' ELSE
      expandedKey(109);
  
  out0_109(110) <= out0_108(110) WHEN out0_16 = '0' ELSE
      expandedKey(110);
  
  out0_109(111) <= out0_108(111) WHEN out0_16 = '0' ELSE
      expandedKey(111);
  
  out0_109(112) <= out0_108(112) WHEN out0_16 = '0' ELSE
      expandedKey(112);
  
  out0_109(113) <= out0_108(113) WHEN out0_16 = '0' ELSE
      expandedKey(113);
  
  out0_109(114) <= out0_108(114) WHEN out0_16 = '0' ELSE
      expandedKey(114);
  
  out0_109(115) <= out0_108(115) WHEN out0_16 = '0' ELSE
      expandedKey(115);
  
  out0_109(116) <= out0_108(116) WHEN out0_16 = '0' ELSE
      expandedKey(116);
  
  out0_109(117) <= out0_108(117) WHEN out0_16 = '0' ELSE
      expandedKey(117);
  
  out0_109(118) <= out0_108(118) WHEN out0_16 = '0' ELSE
      expandedKey(118);
  
  out0_109(119) <= out0_108(119) WHEN out0_16 = '0' ELSE
      expandedKey(119);
  
  out0_109(120) <= out0_108(120) WHEN out0_16 = '0' ELSE
      expandedKey(120);
  
  out0_109(121) <= out0_108(121) WHEN out0_16 = '0' ELSE
      expandedKey(121);
  
  out0_109(122) <= out0_108(122) WHEN out0_16 = '0' ELSE
      expandedKey(122);
  
  out0_109(123) <= out0_108(123) WHEN out0_16 = '0' ELSE
      expandedKey(123);
  
  out0_109(124) <= out0_108(124) WHEN out0_16 = '0' ELSE
      expandedKey(124);
  
  out0_109(125) <= out0_108(125) WHEN out0_16 = '0' ELSE
      expandedKey(125);
  
  out0_109(126) <= out0_108(126) WHEN out0_16 = '0' ELSE
      expandedKey(126);
  
  out0_109(127) <= out0_108(127) WHEN out0_16 = '0' ELSE
      expandedKey(127);
  
  out0_109(128) <= out0_108(128) WHEN out0_16 = '0' ELSE
      expandedKey(128);
  
  out0_109(129) <= out0_108(129) WHEN out0_16 = '0' ELSE
      expandedKey(129);
  
  out0_109(130) <= out0_108(130) WHEN out0_16 = '0' ELSE
      expandedKey(130);
  
  out0_109(131) <= out0_108(131) WHEN out0_16 = '0' ELSE
      expandedKey(131);
  
  out0_109(132) <= out0_108(132) WHEN out0_16 = '0' ELSE
      expandedKey(132);
  
  out0_109(133) <= out0_108(133) WHEN out0_16 = '0' ELSE
      expandedKey(133);
  
  out0_109(134) <= out0_108(134) WHEN out0_16 = '0' ELSE
      expandedKey(134);
  
  out0_109(135) <= out0_108(135) WHEN out0_16 = '0' ELSE
      expandedKey(135);
  
  out0_109(136) <= out0_108(136) WHEN out0_16 = '0' ELSE
      expandedKey(136);
  
  out0_109(137) <= out0_108(137) WHEN out0_16 = '0' ELSE
      expandedKey(137);
  
  out0_109(138) <= out0_108(138) WHEN out0_16 = '0' ELSE
      expandedKey(138);
  
  out0_109(139) <= out0_108(139) WHEN out0_16 = '0' ELSE
      expandedKey(139);
  
  out0_109(140) <= out0_108(140) WHEN out0_16 = '0' ELSE
      expandedKey(140);
  
  out0_109(141) <= out0_108(141) WHEN out0_16 = '0' ELSE
      expandedKey(141);
  
  out0_109(142) <= out0_108(142) WHEN out0_16 = '0' ELSE
      expandedKey(142);
  
  out0_109(143) <= out0_108(143) WHEN out0_16 = '0' ELSE
      expandedKey(143);
  
  out0_109(144) <= out0_108(144) WHEN out0_16 = '0' ELSE
      expandedKey(144);
  
  out0_109(145) <= out0_108(145) WHEN out0_16 = '0' ELSE
      expandedKey(145);
  
  out0_109(146) <= out0_108(146) WHEN out0_16 = '0' ELSE
      expandedKey(146);
  
  out0_109(147) <= out0_108(147) WHEN out0_16 = '0' ELSE
      expandedKey(147);
  
  out0_109(148) <= out0_108(148) WHEN out0_16 = '0' ELSE
      expandedKey(148);
  
  out0_109(149) <= out0_108(149) WHEN out0_16 = '0' ELSE
      expandedKey(149);
  
  out0_109(150) <= out0_108(150) WHEN out0_16 = '0' ELSE
      expandedKey(150);
  
  out0_109(151) <= out0_108(151) WHEN out0_16 = '0' ELSE
      expandedKey(151);
  
  out0_109(152) <= out0_108(152) WHEN out0_16 = '0' ELSE
      expandedKey(152);
  
  out0_109(153) <= out0_108(153) WHEN out0_16 = '0' ELSE
      expandedKey(153);
  
  out0_109(154) <= out0_108(154) WHEN out0_16 = '0' ELSE
      expandedKey(154);
  
  out0_109(155) <= out0_108(155) WHEN out0_16 = '0' ELSE
      expandedKey(155);
  
  out0_109(156) <= out0_108(156) WHEN out0_16 = '0' ELSE
      expandedKey(156);
  
  out0_109(157) <= out0_108(157) WHEN out0_16 = '0' ELSE
      expandedKey(157);
  
  out0_109(158) <= out0_108(158) WHEN out0_16 = '0' ELSE
      expandedKey(158);
  
  out0_109(159) <= out0_108(159) WHEN out0_16 = '0' ELSE
      expandedKey(159);
  
  out0_109(160) <= out0_108(160) WHEN out0_16 = '0' ELSE
      expandedKey(160);
  
  out0_109(161) <= out0_108(161) WHEN out0_16 = '0' ELSE
      expandedKey(161);
  
  out0_109(162) <= out0_108(162) WHEN out0_16 = '0' ELSE
      expandedKey(162);
  
  out0_109(163) <= out0_108(163) WHEN out0_16 = '0' ELSE
      expandedKey(163);
  
  out0_109(164) <= out0_108(164) WHEN out0_16 = '0' ELSE
      expandedKey(164);
  
  out0_109(165) <= out0_108(165) WHEN out0_16 = '0' ELSE
      expandedKey(165);
  
  out0_109(166) <= out0_108(166) WHEN out0_16 = '0' ELSE
      expandedKey(166);
  
  out0_109(167) <= out0_108(167) WHEN out0_16 = '0' ELSE
      expandedKey(167);
  
  out0_109(168) <= out0_108(168) WHEN out0_16 = '0' ELSE
      expandedKey(168);
  
  out0_109(169) <= out0_108(169) WHEN out0_16 = '0' ELSE
      expandedKey(169);
  
  out0_109(170) <= out0_108(170) WHEN out0_16 = '0' ELSE
      expandedKey(170);
  
  out0_109(171) <= out0_108(171) WHEN out0_16 = '0' ELSE
      expandedKey(171);
  
  out0_109(172) <= out0_108(172) WHEN out0_16 = '0' ELSE
      expandedKey(172);
  
  out0_109(173) <= out0_108(173) WHEN out0_16 = '0' ELSE
      expandedKey(173);
  
  out0_109(174) <= out0_108(174) WHEN out0_16 = '0' ELSE
      expandedKey(174);
  
  out0_109(175) <= out0_108(175) WHEN out0_16 = '0' ELSE
      expandedKey(175);
  
  out0_109(176) <= out0_108(176) WHEN out0_16 = '0' ELSE
      expandedKey(176);
  
  out0_109(177) <= out0_108(177) WHEN out0_16 = '0' ELSE
      expandedKey(177);
  
  out0_109(178) <= out0_108(178) WHEN out0_16 = '0' ELSE
      expandedKey(178);
  
  out0_109(179) <= out0_108(179) WHEN out0_16 = '0' ELSE
      expandedKey(179);
  
  out0_109(180) <= out0_108(180) WHEN out0_16 = '0' ELSE
      expandedKey(180);
  
  out0_109(181) <= out0_108(181) WHEN out0_16 = '0' ELSE
      expandedKey(181);
  
  out0_109(182) <= out0_108(182) WHEN out0_16 = '0' ELSE
      expandedKey(182);
  
  out0_109(183) <= out0_108(183) WHEN out0_16 = '0' ELSE
      expandedKey(183);
  
  out0_109(184) <= out0_108(184) WHEN out0_16 = '0' ELSE
      expandedKey(184);
  
  out0_109(185) <= out0_108(185) WHEN out0_16 = '0' ELSE
      expandedKey(185);
  
  out0_109(186) <= out0_108(186) WHEN out0_16 = '0' ELSE
      expandedKey(186);
  
  out0_109(187) <= out0_108(187) WHEN out0_16 = '0' ELSE
      expandedKey(187);
  
  out0_109(188) <= out0_108(188) WHEN out0_16 = '0' ELSE
      expandedKey(188);
  
  out0_109(189) <= out0_108(189) WHEN out0_16 = '0' ELSE
      expandedKey(189);
  
  out0_109(190) <= out0_108(190) WHEN out0_16 = '0' ELSE
      expandedKey(190);
  
  out0_109(191) <= out0_108(191) WHEN out0_16 = '0' ELSE
      expandedKey(191);
  
  out0_109(192) <= out0_108(192) WHEN out0_16 = '0' ELSE
      expandedKey(192);
  
  out0_109(193) <= out0_108(193) WHEN out0_16 = '0' ELSE
      expandedKey(193);
  
  out0_109(194) <= out0_108(194) WHEN out0_16 = '0' ELSE
      expandedKey(194);
  
  out0_109(195) <= out0_108(195) WHEN out0_16 = '0' ELSE
      expandedKey(195);
  
  out0_109(196) <= out0_108(196) WHEN out0_16 = '0' ELSE
      expandedKey(196);
  
  out0_109(197) <= out0_108(197) WHEN out0_16 = '0' ELSE
      expandedKey(197);
  
  out0_109(198) <= out0_108(198) WHEN out0_16 = '0' ELSE
      expandedKey(198);
  
  out0_109(199) <= out0_108(199) WHEN out0_16 = '0' ELSE
      expandedKey(199);
  
  out0_109(200) <= out0_108(200) WHEN out0_16 = '0' ELSE
      expandedKey(200);
  
  out0_109(201) <= out0_108(201) WHEN out0_16 = '0' ELSE
      expandedKey(201);
  
  out0_109(202) <= out0_108(202) WHEN out0_16 = '0' ELSE
      expandedKey(202);
  
  out0_109(203) <= out0_108(203) WHEN out0_16 = '0' ELSE
      expandedKey(203);
  
  out0_109(204) <= out0_108(204) WHEN out0_16 = '0' ELSE
      expandedKey(204);
  
  out0_109(205) <= out0_108(205) WHEN out0_16 = '0' ELSE
      expandedKey(205);
  
  out0_109(206) <= out0_108(206) WHEN out0_16 = '0' ELSE
      expandedKey(206);
  
  out0_109(207) <= out0_108(207) WHEN out0_16 = '0' ELSE
      expandedKey(207);
  
  out0_109(208) <= out0_108(208) WHEN out0_16 = '0' ELSE
      expandedKey(208);
  
  out0_109(209) <= out0_108(209) WHEN out0_16 = '0' ELSE
      expandedKey(209);
  
  out0_109(210) <= out0_108(210) WHEN out0_16 = '0' ELSE
      expandedKey(210);
  
  out0_109(211) <= out0_108(211) WHEN out0_16 = '0' ELSE
      expandedKey(211);
  
  out0_109(212) <= out0_108(212) WHEN out0_16 = '0' ELSE
      expandedKey(212);
  
  out0_109(213) <= out0_108(213) WHEN out0_16 = '0' ELSE
      expandedKey(213);
  
  out0_109(214) <= out0_108(214) WHEN out0_16 = '0' ELSE
      expandedKey(214);
  
  out0_109(215) <= out0_108(215) WHEN out0_16 = '0' ELSE
      expandedKey(215);
  
  out0_109(216) <= out0_108(216) WHEN out0_16 = '0' ELSE
      expandedKey(216);
  
  out0_109(217) <= out0_108(217) WHEN out0_16 = '0' ELSE
      expandedKey(217);
  
  out0_109(218) <= out0_108(218) WHEN out0_16 = '0' ELSE
      expandedKey(218);
  
  out0_109(219) <= out0_108(219) WHEN out0_16 = '0' ELSE
      expandedKey(219);
  
  out0_109(220) <= out0_108(220) WHEN out0_16 = '0' ELSE
      expandedKey(220);
  
  out0_109(221) <= out0_108(221) WHEN out0_16 = '0' ELSE
      expandedKey(221);
  
  out0_109(222) <= out0_108(222) WHEN out0_16 = '0' ELSE
      expandedKey(222);
  
  out0_109(223) <= out0_108(223) WHEN out0_16 = '0' ELSE
      expandedKey(223);
  
  out0_109(224) <= out0_108(224) WHEN out0_16 = '0' ELSE
      expandedKey(224);
  
  out0_109(225) <= out0_108(225) WHEN out0_16 = '0' ELSE
      expandedKey(225);
  
  out0_109(226) <= out0_108(226) WHEN out0_16 = '0' ELSE
      expandedKey(226);
  
  out0_109(227) <= out0_108(227) WHEN out0_16 = '0' ELSE
      expandedKey(227);
  
  out0_109(228) <= out0_108(228) WHEN out0_16 = '0' ELSE
      expandedKey(228);
  
  out0_109(229) <= out0_108(229) WHEN out0_16 = '0' ELSE
      expandedKey(229);
  
  out0_109(230) <= out0_108(230) WHEN out0_16 = '0' ELSE
      expandedKey(230);
  
  out0_109(231) <= out0_108(231) WHEN out0_16 = '0' ELSE
      expandedKey(231);
  
  out0_109(232) <= out0_108(232) WHEN out0_16 = '0' ELSE
      expandedKey(232);
  
  out0_109(233) <= out0_108(233) WHEN out0_16 = '0' ELSE
      expandedKey(233);
  
  out0_109(234) <= out0_108(234) WHEN out0_16 = '0' ELSE
      expandedKey(234);
  
  out0_109(235) <= out0_108(235) WHEN out0_16 = '0' ELSE
      expandedKey(235);
  
  out0_109(236) <= out0_108(236) WHEN out0_16 = '0' ELSE
      expandedKey(236);
  
  out0_109(237) <= out0_108(237) WHEN out0_16 = '0' ELSE
      expandedKey(237);
  
  out0_109(238) <= out0_108(238) WHEN out0_16 = '0' ELSE
      expandedKey(238);
  
  out0_109(239) <= out0_108(239) WHEN out0_16 = '0' ELSE
      expandedKey(239);

  
  out0_110(0) <= out0_109(0) WHEN out0_18 = '0' ELSE
      expandedKey(0);
  
  out0_110(1) <= out0_109(1) WHEN out0_18 = '0' ELSE
      expandedKey(1);
  
  out0_110(2) <= out0_109(2) WHEN out0_18 = '0' ELSE
      expandedKey(2);
  
  out0_110(3) <= out0_109(3) WHEN out0_18 = '0' ELSE
      expandedKey(3);
  
  out0_110(4) <= out0_109(4) WHEN out0_18 = '0' ELSE
      expandedKey(4);
  
  out0_110(5) <= out0_109(5) WHEN out0_18 = '0' ELSE
      expandedKey(5);
  
  out0_110(6) <= out0_109(6) WHEN out0_18 = '0' ELSE
      expandedKey(6);
  
  out0_110(7) <= out0_109(7) WHEN out0_18 = '0' ELSE
      expandedKey(7);
  
  out0_110(8) <= out0_109(8) WHEN out0_18 = '0' ELSE
      expandedKey(8);
  
  out0_110(9) <= out0_109(9) WHEN out0_18 = '0' ELSE
      expandedKey(9);
  
  out0_110(10) <= out0_109(10) WHEN out0_18 = '0' ELSE
      expandedKey(10);
  
  out0_110(11) <= out0_109(11) WHEN out0_18 = '0' ELSE
      expandedKey(11);
  
  out0_110(12) <= out0_109(12) WHEN out0_18 = '0' ELSE
      expandedKey(12);
  
  out0_110(13) <= out0_109(13) WHEN out0_18 = '0' ELSE
      expandedKey(13);
  
  out0_110(14) <= out0_109(14) WHEN out0_18 = '0' ELSE
      expandedKey(14);
  
  out0_110(15) <= out0_109(15) WHEN out0_18 = '0' ELSE
      expandedKey(15);
  
  out0_110(16) <= out0_109(16) WHEN out0_18 = '0' ELSE
      expandedKey(16);
  
  out0_110(17) <= out0_109(17) WHEN out0_18 = '0' ELSE
      expandedKey(17);
  
  out0_110(18) <= out0_109(18) WHEN out0_18 = '0' ELSE
      expandedKey(18);
  
  out0_110(19) <= out0_109(19) WHEN out0_18 = '0' ELSE
      expandedKey(19);
  
  out0_110(20) <= out0_109(20) WHEN out0_18 = '0' ELSE
      expandedKey(20);
  
  out0_110(21) <= out0_109(21) WHEN out0_18 = '0' ELSE
      expandedKey(21);
  
  out0_110(22) <= out0_109(22) WHEN out0_18 = '0' ELSE
      expandedKey(22);
  
  out0_110(23) <= out0_109(23) WHEN out0_18 = '0' ELSE
      expandedKey(23);
  
  out0_110(24) <= out0_109(24) WHEN out0_18 = '0' ELSE
      expandedKey(24);
  
  out0_110(25) <= out0_109(25) WHEN out0_18 = '0' ELSE
      expandedKey(25);
  
  out0_110(26) <= out0_109(26) WHEN out0_18 = '0' ELSE
      expandedKey(26);
  
  out0_110(27) <= out0_109(27) WHEN out0_18 = '0' ELSE
      expandedKey(27);
  
  out0_110(28) <= out0_109(28) WHEN out0_18 = '0' ELSE
      expandedKey(28);
  
  out0_110(29) <= out0_109(29) WHEN out0_18 = '0' ELSE
      expandedKey(29);
  
  out0_110(30) <= out0_109(30) WHEN out0_18 = '0' ELSE
      expandedKey(30);
  
  out0_110(31) <= out0_109(31) WHEN out0_18 = '0' ELSE
      expandedKey(31);
  
  out0_110(32) <= out0_109(32) WHEN out0_18 = '0' ELSE
      expandedKey(32);
  
  out0_110(33) <= out0_109(33) WHEN out0_18 = '0' ELSE
      expandedKey(33);
  
  out0_110(34) <= out0_109(34) WHEN out0_18 = '0' ELSE
      expandedKey(34);
  
  out0_110(35) <= out0_109(35) WHEN out0_18 = '0' ELSE
      expandedKey(35);
  
  out0_110(36) <= out0_109(36) WHEN out0_18 = '0' ELSE
      expandedKey(36);
  
  out0_110(37) <= out0_109(37) WHEN out0_18 = '0' ELSE
      expandedKey(37);
  
  out0_110(38) <= out0_109(38) WHEN out0_18 = '0' ELSE
      expandedKey(38);
  
  out0_110(39) <= out0_109(39) WHEN out0_18 = '0' ELSE
      expandedKey(39);
  
  out0_110(40) <= out0_109(40) WHEN out0_18 = '0' ELSE
      expandedKey(40);
  
  out0_110(41) <= out0_109(41) WHEN out0_18 = '0' ELSE
      expandedKey(41);
  
  out0_110(42) <= out0_109(42) WHEN out0_18 = '0' ELSE
      expandedKey(42);
  
  out0_110(43) <= out0_109(43) WHEN out0_18 = '0' ELSE
      expandedKey(43);
  
  out0_110(44) <= out0_109(44) WHEN out0_18 = '0' ELSE
      expandedKey(44);
  
  out0_110(45) <= out0_109(45) WHEN out0_18 = '0' ELSE
      expandedKey(45);
  
  out0_110(46) <= out0_109(46) WHEN out0_18 = '0' ELSE
      expandedKey(46);
  
  out0_110(47) <= out0_109(47) WHEN out0_18 = '0' ELSE
      expandedKey(47);
  
  out0_110(48) <= out0_109(48) WHEN out0_18 = '0' ELSE
      expandedKey(48);
  
  out0_110(49) <= out0_109(49) WHEN out0_18 = '0' ELSE
      expandedKey(49);
  
  out0_110(50) <= out0_109(50) WHEN out0_18 = '0' ELSE
      expandedKey(50);
  
  out0_110(51) <= out0_109(51) WHEN out0_18 = '0' ELSE
      expandedKey(51);
  
  out0_110(52) <= out0_109(52) WHEN out0_18 = '0' ELSE
      expandedKey(52);
  
  out0_110(53) <= out0_109(53) WHEN out0_18 = '0' ELSE
      expandedKey(53);
  
  out0_110(54) <= out0_109(54) WHEN out0_18 = '0' ELSE
      expandedKey(54);
  
  out0_110(55) <= out0_109(55) WHEN out0_18 = '0' ELSE
      expandedKey(55);
  
  out0_110(56) <= out0_109(56) WHEN out0_18 = '0' ELSE
      expandedKey(56);
  
  out0_110(57) <= out0_109(57) WHEN out0_18 = '0' ELSE
      expandedKey(57);
  
  out0_110(58) <= out0_109(58) WHEN out0_18 = '0' ELSE
      expandedKey(58);
  
  out0_110(59) <= out0_109(59) WHEN out0_18 = '0' ELSE
      expandedKey(59);
  
  out0_110(60) <= out0_109(60) WHEN out0_18 = '0' ELSE
      expandedKey(60);
  
  out0_110(61) <= out0_109(61) WHEN out0_18 = '0' ELSE
      expandedKey(61);
  
  out0_110(62) <= out0_109(62) WHEN out0_18 = '0' ELSE
      expandedKey(62);
  
  out0_110(63) <= out0_109(63) WHEN out0_18 = '0' ELSE
      expandedKey(63);
  
  out0_110(64) <= out0_109(64) WHEN out0_18 = '0' ELSE
      expandedKey(64);
  
  out0_110(65) <= out0_109(65) WHEN out0_18 = '0' ELSE
      expandedKey(65);
  
  out0_110(66) <= out0_109(66) WHEN out0_18 = '0' ELSE
      expandedKey(66);
  
  out0_110(67) <= out0_109(67) WHEN out0_18 = '0' ELSE
      expandedKey(67);
  
  out0_110(68) <= out0_109(68) WHEN out0_18 = '0' ELSE
      expandedKey(68);
  
  out0_110(69) <= out0_109(69) WHEN out0_18 = '0' ELSE
      expandedKey(69);
  
  out0_110(70) <= out0_109(70) WHEN out0_18 = '0' ELSE
      expandedKey(70);
  
  out0_110(71) <= out0_109(71) WHEN out0_18 = '0' ELSE
      expandedKey(71);
  
  out0_110(72) <= out0_109(72) WHEN out0_18 = '0' ELSE
      expandedKey(72);
  
  out0_110(73) <= out0_109(73) WHEN out0_18 = '0' ELSE
      expandedKey(73);
  
  out0_110(74) <= out0_109(74) WHEN out0_18 = '0' ELSE
      expandedKey(74);
  
  out0_110(75) <= out0_109(75) WHEN out0_18 = '0' ELSE
      expandedKey(75);
  
  out0_110(76) <= out0_109(76) WHEN out0_18 = '0' ELSE
      expandedKey(76);
  
  out0_110(77) <= out0_109(77) WHEN out0_18 = '0' ELSE
      expandedKey(77);
  
  out0_110(78) <= out0_109(78) WHEN out0_18 = '0' ELSE
      expandedKey(78);
  
  out0_110(79) <= out0_109(79) WHEN out0_18 = '0' ELSE
      expandedKey(79);
  
  out0_110(80) <= out0_109(80) WHEN out0_18 = '0' ELSE
      expandedKey(80);
  
  out0_110(81) <= out0_109(81) WHEN out0_18 = '0' ELSE
      expandedKey(81);
  
  out0_110(82) <= out0_109(82) WHEN out0_18 = '0' ELSE
      expandedKey(82);
  
  out0_110(83) <= out0_109(83) WHEN out0_18 = '0' ELSE
      expandedKey(83);
  
  out0_110(84) <= out0_109(84) WHEN out0_18 = '0' ELSE
      expandedKey(84);
  
  out0_110(85) <= out0_109(85) WHEN out0_18 = '0' ELSE
      expandedKey(85);
  
  out0_110(86) <= out0_109(86) WHEN out0_18 = '0' ELSE
      expandedKey(86);
  
  out0_110(87) <= out0_109(87) WHEN out0_18 = '0' ELSE
      expandedKey(87);
  
  out0_110(88) <= out0_109(88) WHEN out0_18 = '0' ELSE
      expandedKey(88);
  
  out0_110(89) <= out0_109(89) WHEN out0_18 = '0' ELSE
      expandedKey(89);
  
  out0_110(90) <= out0_109(90) WHEN out0_18 = '0' ELSE
      expandedKey(90);
  
  out0_110(91) <= out0_109(91) WHEN out0_18 = '0' ELSE
      expandedKey(91);
  
  out0_110(92) <= out0_109(92) WHEN out0_18 = '0' ELSE
      expandedKey(92);
  
  out0_110(93) <= out0_109(93) WHEN out0_18 = '0' ELSE
      expandedKey(93);
  
  out0_110(94) <= out0_109(94) WHEN out0_18 = '0' ELSE
      expandedKey(94);
  
  out0_110(95) <= out0_109(95) WHEN out0_18 = '0' ELSE
      expandedKey(95);
  
  out0_110(96) <= out0_109(96) WHEN out0_18 = '0' ELSE
      expandedKey(96);
  
  out0_110(97) <= out0_109(97) WHEN out0_18 = '0' ELSE
      expandedKey(97);
  
  out0_110(98) <= out0_109(98) WHEN out0_18 = '0' ELSE
      expandedKey(98);
  
  out0_110(99) <= out0_109(99) WHEN out0_18 = '0' ELSE
      expandedKey(99);
  
  out0_110(100) <= out0_109(100) WHEN out0_18 = '0' ELSE
      expandedKey(100);
  
  out0_110(101) <= out0_109(101) WHEN out0_18 = '0' ELSE
      expandedKey(101);
  
  out0_110(102) <= out0_109(102) WHEN out0_18 = '0' ELSE
      expandedKey(102);
  
  out0_110(103) <= out0_109(103) WHEN out0_18 = '0' ELSE
      expandedKey(103);
  
  out0_110(104) <= out0_109(104) WHEN out0_18 = '0' ELSE
      expandedKey(104);
  
  out0_110(105) <= out0_109(105) WHEN out0_18 = '0' ELSE
      expandedKey(105);
  
  out0_110(106) <= out0_109(106) WHEN out0_18 = '0' ELSE
      expandedKey(106);
  
  out0_110(107) <= out0_109(107) WHEN out0_18 = '0' ELSE
      expandedKey(107);
  
  out0_110(108) <= out0_109(108) WHEN out0_18 = '0' ELSE
      expandedKey(108);
  
  out0_110(109) <= out0_109(109) WHEN out0_18 = '0' ELSE
      expandedKey(109);
  
  out0_110(110) <= out0_109(110) WHEN out0_18 = '0' ELSE
      expandedKey(110);
  
  out0_110(111) <= out0_109(111) WHEN out0_18 = '0' ELSE
      expandedKey(111);
  
  out0_110(112) <= out0_109(112) WHEN out0_18 = '0' ELSE
      expandedKey(112);
  
  out0_110(113) <= out0_109(113) WHEN out0_18 = '0' ELSE
      expandedKey(113);
  
  out0_110(114) <= out0_109(114) WHEN out0_18 = '0' ELSE
      expandedKey(114);
  
  out0_110(115) <= out0_109(115) WHEN out0_18 = '0' ELSE
      expandedKey(115);
  
  out0_110(116) <= out0_109(116) WHEN out0_18 = '0' ELSE
      expandedKey(116);
  
  out0_110(117) <= out0_109(117) WHEN out0_18 = '0' ELSE
      expandedKey(117);
  
  out0_110(118) <= out0_109(118) WHEN out0_18 = '0' ELSE
      expandedKey(118);
  
  out0_110(119) <= out0_109(119) WHEN out0_18 = '0' ELSE
      expandedKey(119);
  
  out0_110(120) <= out0_109(120) WHEN out0_18 = '0' ELSE
      expandedKey(120);
  
  out0_110(121) <= out0_109(121) WHEN out0_18 = '0' ELSE
      expandedKey(121);
  
  out0_110(122) <= out0_109(122) WHEN out0_18 = '0' ELSE
      expandedKey(122);
  
  out0_110(123) <= out0_109(123) WHEN out0_18 = '0' ELSE
      expandedKey(123);
  
  out0_110(124) <= out0_109(124) WHEN out0_18 = '0' ELSE
      expandedKey(124);
  
  out0_110(125) <= out0_109(125) WHEN out0_18 = '0' ELSE
      expandedKey(125);
  
  out0_110(126) <= out0_109(126) WHEN out0_18 = '0' ELSE
      expandedKey(126);
  
  out0_110(127) <= out0_109(127) WHEN out0_18 = '0' ELSE
      expandedKey(127);
  
  out0_110(128) <= out0_109(128) WHEN out0_18 = '0' ELSE
      expandedKey(128);
  
  out0_110(129) <= out0_109(129) WHEN out0_18 = '0' ELSE
      expandedKey(129);
  
  out0_110(130) <= out0_109(130) WHEN out0_18 = '0' ELSE
      expandedKey(130);
  
  out0_110(131) <= out0_109(131) WHEN out0_18 = '0' ELSE
      expandedKey(131);
  
  out0_110(132) <= out0_109(132) WHEN out0_18 = '0' ELSE
      expandedKey(132);
  
  out0_110(133) <= out0_109(133) WHEN out0_18 = '0' ELSE
      expandedKey(133);
  
  out0_110(134) <= out0_109(134) WHEN out0_18 = '0' ELSE
      expandedKey(134);
  
  out0_110(135) <= out0_109(135) WHEN out0_18 = '0' ELSE
      expandedKey(135);
  
  out0_110(136) <= out0_109(136) WHEN out0_18 = '0' ELSE
      expandedKey(136);
  
  out0_110(137) <= out0_109(137) WHEN out0_18 = '0' ELSE
      expandedKey(137);
  
  out0_110(138) <= out0_109(138) WHEN out0_18 = '0' ELSE
      expandedKey(138);
  
  out0_110(139) <= out0_109(139) WHEN out0_18 = '0' ELSE
      expandedKey(139);
  
  out0_110(140) <= out0_109(140) WHEN out0_18 = '0' ELSE
      expandedKey(140);
  
  out0_110(141) <= out0_109(141) WHEN out0_18 = '0' ELSE
      expandedKey(141);
  
  out0_110(142) <= out0_109(142) WHEN out0_18 = '0' ELSE
      expandedKey(142);
  
  out0_110(143) <= out0_109(143) WHEN out0_18 = '0' ELSE
      expandedKey(143);
  
  out0_110(144) <= out0_109(144) WHEN out0_18 = '0' ELSE
      expandedKey(144);
  
  out0_110(145) <= out0_109(145) WHEN out0_18 = '0' ELSE
      expandedKey(145);
  
  out0_110(146) <= out0_109(146) WHEN out0_18 = '0' ELSE
      expandedKey(146);
  
  out0_110(147) <= out0_109(147) WHEN out0_18 = '0' ELSE
      expandedKey(147);
  
  out0_110(148) <= out0_109(148) WHEN out0_18 = '0' ELSE
      expandedKey(148);
  
  out0_110(149) <= out0_109(149) WHEN out0_18 = '0' ELSE
      expandedKey(149);
  
  out0_110(150) <= out0_109(150) WHEN out0_18 = '0' ELSE
      expandedKey(150);
  
  out0_110(151) <= out0_109(151) WHEN out0_18 = '0' ELSE
      expandedKey(151);
  
  out0_110(152) <= out0_109(152) WHEN out0_18 = '0' ELSE
      expandedKey(152);
  
  out0_110(153) <= out0_109(153) WHEN out0_18 = '0' ELSE
      expandedKey(153);
  
  out0_110(154) <= out0_109(154) WHEN out0_18 = '0' ELSE
      expandedKey(154);
  
  out0_110(155) <= out0_109(155) WHEN out0_18 = '0' ELSE
      expandedKey(155);
  
  out0_110(156) <= out0_109(156) WHEN out0_18 = '0' ELSE
      expandedKey(156);
  
  out0_110(157) <= out0_109(157) WHEN out0_18 = '0' ELSE
      expandedKey(157);
  
  out0_110(158) <= out0_109(158) WHEN out0_18 = '0' ELSE
      expandedKey(158);
  
  out0_110(159) <= out0_109(159) WHEN out0_18 = '0' ELSE
      expandedKey(159);
  
  out0_110(160) <= out0_109(160) WHEN out0_18 = '0' ELSE
      expandedKey(160);
  
  out0_110(161) <= out0_109(161) WHEN out0_18 = '0' ELSE
      expandedKey(161);
  
  out0_110(162) <= out0_109(162) WHEN out0_18 = '0' ELSE
      expandedKey(162);
  
  out0_110(163) <= out0_109(163) WHEN out0_18 = '0' ELSE
      expandedKey(163);
  
  out0_110(164) <= out0_109(164) WHEN out0_18 = '0' ELSE
      expandedKey(164);
  
  out0_110(165) <= out0_109(165) WHEN out0_18 = '0' ELSE
      expandedKey(165);
  
  out0_110(166) <= out0_109(166) WHEN out0_18 = '0' ELSE
      expandedKey(166);
  
  out0_110(167) <= out0_109(167) WHEN out0_18 = '0' ELSE
      expandedKey(167);
  
  out0_110(168) <= out0_109(168) WHEN out0_18 = '0' ELSE
      expandedKey(168);
  
  out0_110(169) <= out0_109(169) WHEN out0_18 = '0' ELSE
      expandedKey(169);
  
  out0_110(170) <= out0_109(170) WHEN out0_18 = '0' ELSE
      expandedKey(170);
  
  out0_110(171) <= out0_109(171) WHEN out0_18 = '0' ELSE
      expandedKey(171);
  
  out0_110(172) <= out0_109(172) WHEN out0_18 = '0' ELSE
      expandedKey(172);
  
  out0_110(173) <= out0_109(173) WHEN out0_18 = '0' ELSE
      expandedKey(173);
  
  out0_110(174) <= out0_109(174) WHEN out0_18 = '0' ELSE
      expandedKey(174);
  
  out0_110(175) <= out0_109(175) WHEN out0_18 = '0' ELSE
      expandedKey(175);
  
  out0_110(176) <= out0_109(176) WHEN out0_18 = '0' ELSE
      expandedKey(176);
  
  out0_110(177) <= out0_109(177) WHEN out0_18 = '0' ELSE
      expandedKey(177);
  
  out0_110(178) <= out0_109(178) WHEN out0_18 = '0' ELSE
      expandedKey(178);
  
  out0_110(179) <= out0_109(179) WHEN out0_18 = '0' ELSE
      expandedKey(179);
  
  out0_110(180) <= out0_109(180) WHEN out0_18 = '0' ELSE
      expandedKey(180);
  
  out0_110(181) <= out0_109(181) WHEN out0_18 = '0' ELSE
      expandedKey(181);
  
  out0_110(182) <= out0_109(182) WHEN out0_18 = '0' ELSE
      expandedKey(182);
  
  out0_110(183) <= out0_109(183) WHEN out0_18 = '0' ELSE
      expandedKey(183);
  
  out0_110(184) <= out0_109(184) WHEN out0_18 = '0' ELSE
      expandedKey(184);
  
  out0_110(185) <= out0_109(185) WHEN out0_18 = '0' ELSE
      expandedKey(185);
  
  out0_110(186) <= out0_109(186) WHEN out0_18 = '0' ELSE
      expandedKey(186);
  
  out0_110(187) <= out0_109(187) WHEN out0_18 = '0' ELSE
      expandedKey(187);
  
  out0_110(188) <= out0_109(188) WHEN out0_18 = '0' ELSE
      expandedKey(188);
  
  out0_110(189) <= out0_109(189) WHEN out0_18 = '0' ELSE
      expandedKey(189);
  
  out0_110(190) <= out0_109(190) WHEN out0_18 = '0' ELSE
      expandedKey(190);
  
  out0_110(191) <= out0_109(191) WHEN out0_18 = '0' ELSE
      expandedKey(191);
  
  out0_110(192) <= out0_109(192) WHEN out0_18 = '0' ELSE
      expandedKey(192);
  
  out0_110(193) <= out0_109(193) WHEN out0_18 = '0' ELSE
      expandedKey(193);
  
  out0_110(194) <= out0_109(194) WHEN out0_18 = '0' ELSE
      expandedKey(194);
  
  out0_110(195) <= out0_109(195) WHEN out0_18 = '0' ELSE
      expandedKey(195);
  
  out0_110(196) <= out0_109(196) WHEN out0_18 = '0' ELSE
      expandedKey(196);
  
  out0_110(197) <= out0_109(197) WHEN out0_18 = '0' ELSE
      expandedKey(197);
  
  out0_110(198) <= out0_109(198) WHEN out0_18 = '0' ELSE
      expandedKey(198);
  
  out0_110(199) <= out0_109(199) WHEN out0_18 = '0' ELSE
      expandedKey(199);
  
  out0_110(200) <= out0_109(200) WHEN out0_18 = '0' ELSE
      expandedKey(200);
  
  out0_110(201) <= out0_109(201) WHEN out0_18 = '0' ELSE
      expandedKey(201);
  
  out0_110(202) <= out0_109(202) WHEN out0_18 = '0' ELSE
      expandedKey(202);
  
  out0_110(203) <= out0_109(203) WHEN out0_18 = '0' ELSE
      expandedKey(203);
  
  out0_110(204) <= out0_109(204) WHEN out0_18 = '0' ELSE
      expandedKey(204);
  
  out0_110(205) <= out0_109(205) WHEN out0_18 = '0' ELSE
      expandedKey(205);
  
  out0_110(206) <= out0_109(206) WHEN out0_18 = '0' ELSE
      expandedKey(206);
  
  out0_110(207) <= out0_109(207) WHEN out0_18 = '0' ELSE
      expandedKey(207);
  
  out0_110(208) <= out0_109(208) WHEN out0_18 = '0' ELSE
      expandedKey(208);
  
  out0_110(209) <= out0_109(209) WHEN out0_18 = '0' ELSE
      expandedKey(209);
  
  out0_110(210) <= out0_109(210) WHEN out0_18 = '0' ELSE
      expandedKey(210);
  
  out0_110(211) <= out0_109(211) WHEN out0_18 = '0' ELSE
      expandedKey(211);
  
  out0_110(212) <= out0_109(212) WHEN out0_18 = '0' ELSE
      expandedKey(212);
  
  out0_110(213) <= out0_109(213) WHEN out0_18 = '0' ELSE
      expandedKey(213);
  
  out0_110(214) <= out0_109(214) WHEN out0_18 = '0' ELSE
      expandedKey(214);
  
  out0_110(215) <= out0_109(215) WHEN out0_18 = '0' ELSE
      expandedKey(215);
  
  out0_110(216) <= out0_109(216) WHEN out0_18 = '0' ELSE
      expandedKey(216);
  
  out0_110(217) <= out0_109(217) WHEN out0_18 = '0' ELSE
      expandedKey(217);
  
  out0_110(218) <= out0_109(218) WHEN out0_18 = '0' ELSE
      expandedKey(218);
  
  out0_110(219) <= out0_109(219) WHEN out0_18 = '0' ELSE
      expandedKey(219);
  
  out0_110(220) <= out0_109(220) WHEN out0_18 = '0' ELSE
      expandedKey(220);
  
  out0_110(221) <= out0_109(221) WHEN out0_18 = '0' ELSE
      expandedKey(221);
  
  out0_110(222) <= out0_109(222) WHEN out0_18 = '0' ELSE
      expandedKey(222);
  
  out0_110(223) <= out0_109(223) WHEN out0_18 = '0' ELSE
      expandedKey(223);
  
  out0_110(224) <= out0_109(224) WHEN out0_18 = '0' ELSE
      expandedKey(224);
  
  out0_110(225) <= out0_109(225) WHEN out0_18 = '0' ELSE
      expandedKey(225);
  
  out0_110(226) <= out0_109(226) WHEN out0_18 = '0' ELSE
      expandedKey(226);
  
  out0_110(227) <= out0_109(227) WHEN out0_18 = '0' ELSE
      expandedKey(227);
  
  out0_110(228) <= out0_109(228) WHEN out0_18 = '0' ELSE
      expandedKey(228);
  
  out0_110(229) <= out0_109(229) WHEN out0_18 = '0' ELSE
      expandedKey(229);
  
  out0_110(230) <= out0_109(230) WHEN out0_18 = '0' ELSE
      expandedKey(230);
  
  out0_110(231) <= out0_109(231) WHEN out0_18 = '0' ELSE
      expandedKey(231);
  
  out0_110(232) <= out0_109(232) WHEN out0_18 = '0' ELSE
      expandedKey(232);
  
  out0_110(233) <= out0_109(233) WHEN out0_18 = '0' ELSE
      expandedKey(233);
  
  out0_110(234) <= out0_109(234) WHEN out0_18 = '0' ELSE
      expandedKey(234);
  
  out0_110(235) <= out0_109(235) WHEN out0_18 = '0' ELSE
      expandedKey(235);
  
  out0_110(236) <= out0_109(236) WHEN out0_18 = '0' ELSE
      expandedKey(236);
  
  out0_110(237) <= out0_109(237) WHEN out0_18 = '0' ELSE
      expandedKey(237);
  
  out0_110(238) <= out0_109(238) WHEN out0_18 = '0' ELSE
      expandedKey(238);
  
  out0_110(239) <= out0_109(239) WHEN out0_18 = '0' ELSE
      expandedKey(239);

  
  out0_111(0) <= out0_110(0) WHEN out0_20 = '0' ELSE
      expandedKey(0);
  
  out0_111(1) <= out0_110(1) WHEN out0_20 = '0' ELSE
      expandedKey(1);
  
  out0_111(2) <= out0_110(2) WHEN out0_20 = '0' ELSE
      expandedKey(2);
  
  out0_111(3) <= out0_110(3) WHEN out0_20 = '0' ELSE
      expandedKey(3);
  
  out0_111(4) <= out0_110(4) WHEN out0_20 = '0' ELSE
      expandedKey(4);
  
  out0_111(5) <= out0_110(5) WHEN out0_20 = '0' ELSE
      expandedKey(5);
  
  out0_111(6) <= out0_110(6) WHEN out0_20 = '0' ELSE
      expandedKey(6);
  
  out0_111(7) <= out0_110(7) WHEN out0_20 = '0' ELSE
      expandedKey(7);
  
  out0_111(8) <= out0_110(8) WHEN out0_20 = '0' ELSE
      expandedKey(8);
  
  out0_111(9) <= out0_110(9) WHEN out0_20 = '0' ELSE
      expandedKey(9);
  
  out0_111(10) <= out0_110(10) WHEN out0_20 = '0' ELSE
      expandedKey(10);
  
  out0_111(11) <= out0_110(11) WHEN out0_20 = '0' ELSE
      expandedKey(11);
  
  out0_111(12) <= out0_110(12) WHEN out0_20 = '0' ELSE
      expandedKey(12);
  
  out0_111(13) <= out0_110(13) WHEN out0_20 = '0' ELSE
      expandedKey(13);
  
  out0_111(14) <= out0_110(14) WHEN out0_20 = '0' ELSE
      expandedKey(14);
  
  out0_111(15) <= out0_110(15) WHEN out0_20 = '0' ELSE
      expandedKey(15);
  
  out0_111(16) <= out0_110(16) WHEN out0_20 = '0' ELSE
      expandedKey(16);
  
  out0_111(17) <= out0_110(17) WHEN out0_20 = '0' ELSE
      expandedKey(17);
  
  out0_111(18) <= out0_110(18) WHEN out0_20 = '0' ELSE
      expandedKey(18);
  
  out0_111(19) <= out0_110(19) WHEN out0_20 = '0' ELSE
      expandedKey(19);
  
  out0_111(20) <= out0_110(20) WHEN out0_20 = '0' ELSE
      expandedKey(20);
  
  out0_111(21) <= out0_110(21) WHEN out0_20 = '0' ELSE
      expandedKey(21);
  
  out0_111(22) <= out0_110(22) WHEN out0_20 = '0' ELSE
      expandedKey(22);
  
  out0_111(23) <= out0_110(23) WHEN out0_20 = '0' ELSE
      expandedKey(23);
  
  out0_111(24) <= out0_110(24) WHEN out0_20 = '0' ELSE
      expandedKey(24);
  
  out0_111(25) <= out0_110(25) WHEN out0_20 = '0' ELSE
      expandedKey(25);
  
  out0_111(26) <= out0_110(26) WHEN out0_20 = '0' ELSE
      expandedKey(26);
  
  out0_111(27) <= out0_110(27) WHEN out0_20 = '0' ELSE
      expandedKey(27);
  
  out0_111(28) <= out0_110(28) WHEN out0_20 = '0' ELSE
      expandedKey(28);
  
  out0_111(29) <= out0_110(29) WHEN out0_20 = '0' ELSE
      expandedKey(29);
  
  out0_111(30) <= out0_110(30) WHEN out0_20 = '0' ELSE
      expandedKey(30);
  
  out0_111(31) <= out0_110(31) WHEN out0_20 = '0' ELSE
      expandedKey(31);
  
  out0_111(32) <= out0_110(32) WHEN out0_20 = '0' ELSE
      expandedKey(32);
  
  out0_111(33) <= out0_110(33) WHEN out0_20 = '0' ELSE
      expandedKey(33);
  
  out0_111(34) <= out0_110(34) WHEN out0_20 = '0' ELSE
      expandedKey(34);
  
  out0_111(35) <= out0_110(35) WHEN out0_20 = '0' ELSE
      expandedKey(35);
  
  out0_111(36) <= out0_110(36) WHEN out0_20 = '0' ELSE
      expandedKey(36);
  
  out0_111(37) <= out0_110(37) WHEN out0_20 = '0' ELSE
      expandedKey(37);
  
  out0_111(38) <= out0_110(38) WHEN out0_20 = '0' ELSE
      expandedKey(38);
  
  out0_111(39) <= out0_110(39) WHEN out0_20 = '0' ELSE
      expandedKey(39);
  
  out0_111(40) <= out0_110(40) WHEN out0_20 = '0' ELSE
      expandedKey(40);
  
  out0_111(41) <= out0_110(41) WHEN out0_20 = '0' ELSE
      expandedKey(41);
  
  out0_111(42) <= out0_110(42) WHEN out0_20 = '0' ELSE
      expandedKey(42);
  
  out0_111(43) <= out0_110(43) WHEN out0_20 = '0' ELSE
      expandedKey(43);
  
  out0_111(44) <= out0_110(44) WHEN out0_20 = '0' ELSE
      expandedKey(44);
  
  out0_111(45) <= out0_110(45) WHEN out0_20 = '0' ELSE
      expandedKey(45);
  
  out0_111(46) <= out0_110(46) WHEN out0_20 = '0' ELSE
      expandedKey(46);
  
  out0_111(47) <= out0_110(47) WHEN out0_20 = '0' ELSE
      expandedKey(47);
  
  out0_111(48) <= out0_110(48) WHEN out0_20 = '0' ELSE
      expandedKey(48);
  
  out0_111(49) <= out0_110(49) WHEN out0_20 = '0' ELSE
      expandedKey(49);
  
  out0_111(50) <= out0_110(50) WHEN out0_20 = '0' ELSE
      expandedKey(50);
  
  out0_111(51) <= out0_110(51) WHEN out0_20 = '0' ELSE
      expandedKey(51);
  
  out0_111(52) <= out0_110(52) WHEN out0_20 = '0' ELSE
      expandedKey(52);
  
  out0_111(53) <= out0_110(53) WHEN out0_20 = '0' ELSE
      expandedKey(53);
  
  out0_111(54) <= out0_110(54) WHEN out0_20 = '0' ELSE
      expandedKey(54);
  
  out0_111(55) <= out0_110(55) WHEN out0_20 = '0' ELSE
      expandedKey(55);
  
  out0_111(56) <= out0_110(56) WHEN out0_20 = '0' ELSE
      expandedKey(56);
  
  out0_111(57) <= out0_110(57) WHEN out0_20 = '0' ELSE
      expandedKey(57);
  
  out0_111(58) <= out0_110(58) WHEN out0_20 = '0' ELSE
      expandedKey(58);
  
  out0_111(59) <= out0_110(59) WHEN out0_20 = '0' ELSE
      expandedKey(59);
  
  out0_111(60) <= out0_110(60) WHEN out0_20 = '0' ELSE
      expandedKey(60);
  
  out0_111(61) <= out0_110(61) WHEN out0_20 = '0' ELSE
      expandedKey(61);
  
  out0_111(62) <= out0_110(62) WHEN out0_20 = '0' ELSE
      expandedKey(62);
  
  out0_111(63) <= out0_110(63) WHEN out0_20 = '0' ELSE
      expandedKey(63);
  
  out0_111(64) <= out0_110(64) WHEN out0_20 = '0' ELSE
      expandedKey(64);
  
  out0_111(65) <= out0_110(65) WHEN out0_20 = '0' ELSE
      expandedKey(65);
  
  out0_111(66) <= out0_110(66) WHEN out0_20 = '0' ELSE
      expandedKey(66);
  
  out0_111(67) <= out0_110(67) WHEN out0_20 = '0' ELSE
      expandedKey(67);
  
  out0_111(68) <= out0_110(68) WHEN out0_20 = '0' ELSE
      expandedKey(68);
  
  out0_111(69) <= out0_110(69) WHEN out0_20 = '0' ELSE
      expandedKey(69);
  
  out0_111(70) <= out0_110(70) WHEN out0_20 = '0' ELSE
      expandedKey(70);
  
  out0_111(71) <= out0_110(71) WHEN out0_20 = '0' ELSE
      expandedKey(71);
  
  out0_111(72) <= out0_110(72) WHEN out0_20 = '0' ELSE
      expandedKey(72);
  
  out0_111(73) <= out0_110(73) WHEN out0_20 = '0' ELSE
      expandedKey(73);
  
  out0_111(74) <= out0_110(74) WHEN out0_20 = '0' ELSE
      expandedKey(74);
  
  out0_111(75) <= out0_110(75) WHEN out0_20 = '0' ELSE
      expandedKey(75);
  
  out0_111(76) <= out0_110(76) WHEN out0_20 = '0' ELSE
      expandedKey(76);
  
  out0_111(77) <= out0_110(77) WHEN out0_20 = '0' ELSE
      expandedKey(77);
  
  out0_111(78) <= out0_110(78) WHEN out0_20 = '0' ELSE
      expandedKey(78);
  
  out0_111(79) <= out0_110(79) WHEN out0_20 = '0' ELSE
      expandedKey(79);
  
  out0_111(80) <= out0_110(80) WHEN out0_20 = '0' ELSE
      expandedKey(80);
  
  out0_111(81) <= out0_110(81) WHEN out0_20 = '0' ELSE
      expandedKey(81);
  
  out0_111(82) <= out0_110(82) WHEN out0_20 = '0' ELSE
      expandedKey(82);
  
  out0_111(83) <= out0_110(83) WHEN out0_20 = '0' ELSE
      expandedKey(83);
  
  out0_111(84) <= out0_110(84) WHEN out0_20 = '0' ELSE
      expandedKey(84);
  
  out0_111(85) <= out0_110(85) WHEN out0_20 = '0' ELSE
      expandedKey(85);
  
  out0_111(86) <= out0_110(86) WHEN out0_20 = '0' ELSE
      expandedKey(86);
  
  out0_111(87) <= out0_110(87) WHEN out0_20 = '0' ELSE
      expandedKey(87);
  
  out0_111(88) <= out0_110(88) WHEN out0_20 = '0' ELSE
      expandedKey(88);
  
  out0_111(89) <= out0_110(89) WHEN out0_20 = '0' ELSE
      expandedKey(89);
  
  out0_111(90) <= out0_110(90) WHEN out0_20 = '0' ELSE
      expandedKey(90);
  
  out0_111(91) <= out0_110(91) WHEN out0_20 = '0' ELSE
      expandedKey(91);
  
  out0_111(92) <= out0_110(92) WHEN out0_20 = '0' ELSE
      expandedKey(92);
  
  out0_111(93) <= out0_110(93) WHEN out0_20 = '0' ELSE
      expandedKey(93);
  
  out0_111(94) <= out0_110(94) WHEN out0_20 = '0' ELSE
      expandedKey(94);
  
  out0_111(95) <= out0_110(95) WHEN out0_20 = '0' ELSE
      expandedKey(95);
  
  out0_111(96) <= out0_110(96) WHEN out0_20 = '0' ELSE
      expandedKey(96);
  
  out0_111(97) <= out0_110(97) WHEN out0_20 = '0' ELSE
      expandedKey(97);
  
  out0_111(98) <= out0_110(98) WHEN out0_20 = '0' ELSE
      expandedKey(98);
  
  out0_111(99) <= out0_110(99) WHEN out0_20 = '0' ELSE
      expandedKey(99);
  
  out0_111(100) <= out0_110(100) WHEN out0_20 = '0' ELSE
      expandedKey(100);
  
  out0_111(101) <= out0_110(101) WHEN out0_20 = '0' ELSE
      expandedKey(101);
  
  out0_111(102) <= out0_110(102) WHEN out0_20 = '0' ELSE
      expandedKey(102);
  
  out0_111(103) <= out0_110(103) WHEN out0_20 = '0' ELSE
      expandedKey(103);
  
  out0_111(104) <= out0_110(104) WHEN out0_20 = '0' ELSE
      expandedKey(104);
  
  out0_111(105) <= out0_110(105) WHEN out0_20 = '0' ELSE
      expandedKey(105);
  
  out0_111(106) <= out0_110(106) WHEN out0_20 = '0' ELSE
      expandedKey(106);
  
  out0_111(107) <= out0_110(107) WHEN out0_20 = '0' ELSE
      expandedKey(107);
  
  out0_111(108) <= out0_110(108) WHEN out0_20 = '0' ELSE
      expandedKey(108);
  
  out0_111(109) <= out0_110(109) WHEN out0_20 = '0' ELSE
      expandedKey(109);
  
  out0_111(110) <= out0_110(110) WHEN out0_20 = '0' ELSE
      expandedKey(110);
  
  out0_111(111) <= out0_110(111) WHEN out0_20 = '0' ELSE
      expandedKey(111);
  
  out0_111(112) <= out0_110(112) WHEN out0_20 = '0' ELSE
      expandedKey(112);
  
  out0_111(113) <= out0_110(113) WHEN out0_20 = '0' ELSE
      expandedKey(113);
  
  out0_111(114) <= out0_110(114) WHEN out0_20 = '0' ELSE
      expandedKey(114);
  
  out0_111(115) <= out0_110(115) WHEN out0_20 = '0' ELSE
      expandedKey(115);
  
  out0_111(116) <= out0_110(116) WHEN out0_20 = '0' ELSE
      expandedKey(116);
  
  out0_111(117) <= out0_110(117) WHEN out0_20 = '0' ELSE
      expandedKey(117);
  
  out0_111(118) <= out0_110(118) WHEN out0_20 = '0' ELSE
      expandedKey(118);
  
  out0_111(119) <= out0_110(119) WHEN out0_20 = '0' ELSE
      expandedKey(119);
  
  out0_111(120) <= out0_110(120) WHEN out0_20 = '0' ELSE
      expandedKey(120);
  
  out0_111(121) <= out0_110(121) WHEN out0_20 = '0' ELSE
      expandedKey(121);
  
  out0_111(122) <= out0_110(122) WHEN out0_20 = '0' ELSE
      expandedKey(122);
  
  out0_111(123) <= out0_110(123) WHEN out0_20 = '0' ELSE
      expandedKey(123);
  
  out0_111(124) <= out0_110(124) WHEN out0_20 = '0' ELSE
      expandedKey(124);
  
  out0_111(125) <= out0_110(125) WHEN out0_20 = '0' ELSE
      expandedKey(125);
  
  out0_111(126) <= out0_110(126) WHEN out0_20 = '0' ELSE
      expandedKey(126);
  
  out0_111(127) <= out0_110(127) WHEN out0_20 = '0' ELSE
      expandedKey(127);
  
  out0_111(128) <= out0_110(128) WHEN out0_20 = '0' ELSE
      expandedKey(128);
  
  out0_111(129) <= out0_110(129) WHEN out0_20 = '0' ELSE
      expandedKey(129);
  
  out0_111(130) <= out0_110(130) WHEN out0_20 = '0' ELSE
      expandedKey(130);
  
  out0_111(131) <= out0_110(131) WHEN out0_20 = '0' ELSE
      expandedKey(131);
  
  out0_111(132) <= out0_110(132) WHEN out0_20 = '0' ELSE
      expandedKey(132);
  
  out0_111(133) <= out0_110(133) WHEN out0_20 = '0' ELSE
      expandedKey(133);
  
  out0_111(134) <= out0_110(134) WHEN out0_20 = '0' ELSE
      expandedKey(134);
  
  out0_111(135) <= out0_110(135) WHEN out0_20 = '0' ELSE
      expandedKey(135);
  
  out0_111(136) <= out0_110(136) WHEN out0_20 = '0' ELSE
      expandedKey(136);
  
  out0_111(137) <= out0_110(137) WHEN out0_20 = '0' ELSE
      expandedKey(137);
  
  out0_111(138) <= out0_110(138) WHEN out0_20 = '0' ELSE
      expandedKey(138);
  
  out0_111(139) <= out0_110(139) WHEN out0_20 = '0' ELSE
      expandedKey(139);
  
  out0_111(140) <= out0_110(140) WHEN out0_20 = '0' ELSE
      expandedKey(140);
  
  out0_111(141) <= out0_110(141) WHEN out0_20 = '0' ELSE
      expandedKey(141);
  
  out0_111(142) <= out0_110(142) WHEN out0_20 = '0' ELSE
      expandedKey(142);
  
  out0_111(143) <= out0_110(143) WHEN out0_20 = '0' ELSE
      expandedKey(143);
  
  out0_111(144) <= out0_110(144) WHEN out0_20 = '0' ELSE
      expandedKey(144);
  
  out0_111(145) <= out0_110(145) WHEN out0_20 = '0' ELSE
      expandedKey(145);
  
  out0_111(146) <= out0_110(146) WHEN out0_20 = '0' ELSE
      expandedKey(146);
  
  out0_111(147) <= out0_110(147) WHEN out0_20 = '0' ELSE
      expandedKey(147);
  
  out0_111(148) <= out0_110(148) WHEN out0_20 = '0' ELSE
      expandedKey(148);
  
  out0_111(149) <= out0_110(149) WHEN out0_20 = '0' ELSE
      expandedKey(149);
  
  out0_111(150) <= out0_110(150) WHEN out0_20 = '0' ELSE
      expandedKey(150);
  
  out0_111(151) <= out0_110(151) WHEN out0_20 = '0' ELSE
      expandedKey(151);
  
  out0_111(152) <= out0_110(152) WHEN out0_20 = '0' ELSE
      expandedKey(152);
  
  out0_111(153) <= out0_110(153) WHEN out0_20 = '0' ELSE
      expandedKey(153);
  
  out0_111(154) <= out0_110(154) WHEN out0_20 = '0' ELSE
      expandedKey(154);
  
  out0_111(155) <= out0_110(155) WHEN out0_20 = '0' ELSE
      expandedKey(155);
  
  out0_111(156) <= out0_110(156) WHEN out0_20 = '0' ELSE
      expandedKey(156);
  
  out0_111(157) <= out0_110(157) WHEN out0_20 = '0' ELSE
      expandedKey(157);
  
  out0_111(158) <= out0_110(158) WHEN out0_20 = '0' ELSE
      expandedKey(158);
  
  out0_111(159) <= out0_110(159) WHEN out0_20 = '0' ELSE
      expandedKey(159);
  
  out0_111(160) <= out0_110(160) WHEN out0_20 = '0' ELSE
      expandedKey(160);
  
  out0_111(161) <= out0_110(161) WHEN out0_20 = '0' ELSE
      expandedKey(161);
  
  out0_111(162) <= out0_110(162) WHEN out0_20 = '0' ELSE
      expandedKey(162);
  
  out0_111(163) <= out0_110(163) WHEN out0_20 = '0' ELSE
      expandedKey(163);
  
  out0_111(164) <= out0_110(164) WHEN out0_20 = '0' ELSE
      expandedKey(164);
  
  out0_111(165) <= out0_110(165) WHEN out0_20 = '0' ELSE
      expandedKey(165);
  
  out0_111(166) <= out0_110(166) WHEN out0_20 = '0' ELSE
      expandedKey(166);
  
  out0_111(167) <= out0_110(167) WHEN out0_20 = '0' ELSE
      expandedKey(167);
  
  out0_111(168) <= out0_110(168) WHEN out0_20 = '0' ELSE
      expandedKey(168);
  
  out0_111(169) <= out0_110(169) WHEN out0_20 = '0' ELSE
      expandedKey(169);
  
  out0_111(170) <= out0_110(170) WHEN out0_20 = '0' ELSE
      expandedKey(170);
  
  out0_111(171) <= out0_110(171) WHEN out0_20 = '0' ELSE
      expandedKey(171);
  
  out0_111(172) <= out0_110(172) WHEN out0_20 = '0' ELSE
      expandedKey(172);
  
  out0_111(173) <= out0_110(173) WHEN out0_20 = '0' ELSE
      expandedKey(173);
  
  out0_111(174) <= out0_110(174) WHEN out0_20 = '0' ELSE
      expandedKey(174);
  
  out0_111(175) <= out0_110(175) WHEN out0_20 = '0' ELSE
      expandedKey(175);
  
  out0_111(176) <= out0_110(176) WHEN out0_20 = '0' ELSE
      expandedKey(176);
  
  out0_111(177) <= out0_110(177) WHEN out0_20 = '0' ELSE
      expandedKey(177);
  
  out0_111(178) <= out0_110(178) WHEN out0_20 = '0' ELSE
      expandedKey(178);
  
  out0_111(179) <= out0_110(179) WHEN out0_20 = '0' ELSE
      expandedKey(179);
  
  out0_111(180) <= out0_110(180) WHEN out0_20 = '0' ELSE
      expandedKey(180);
  
  out0_111(181) <= out0_110(181) WHEN out0_20 = '0' ELSE
      expandedKey(181);
  
  out0_111(182) <= out0_110(182) WHEN out0_20 = '0' ELSE
      expandedKey(182);
  
  out0_111(183) <= out0_110(183) WHEN out0_20 = '0' ELSE
      expandedKey(183);
  
  out0_111(184) <= out0_110(184) WHEN out0_20 = '0' ELSE
      expandedKey(184);
  
  out0_111(185) <= out0_110(185) WHEN out0_20 = '0' ELSE
      expandedKey(185);
  
  out0_111(186) <= out0_110(186) WHEN out0_20 = '0' ELSE
      expandedKey(186);
  
  out0_111(187) <= out0_110(187) WHEN out0_20 = '0' ELSE
      expandedKey(187);
  
  out0_111(188) <= out0_110(188) WHEN out0_20 = '0' ELSE
      expandedKey(188);
  
  out0_111(189) <= out0_110(189) WHEN out0_20 = '0' ELSE
      expandedKey(189);
  
  out0_111(190) <= out0_110(190) WHEN out0_20 = '0' ELSE
      expandedKey(190);
  
  out0_111(191) <= out0_110(191) WHEN out0_20 = '0' ELSE
      expandedKey(191);
  
  out0_111(192) <= out0_110(192) WHEN out0_20 = '0' ELSE
      expandedKey(192);
  
  out0_111(193) <= out0_110(193) WHEN out0_20 = '0' ELSE
      expandedKey(193);
  
  out0_111(194) <= out0_110(194) WHEN out0_20 = '0' ELSE
      expandedKey(194);
  
  out0_111(195) <= out0_110(195) WHEN out0_20 = '0' ELSE
      expandedKey(195);
  
  out0_111(196) <= out0_110(196) WHEN out0_20 = '0' ELSE
      expandedKey(196);
  
  out0_111(197) <= out0_110(197) WHEN out0_20 = '0' ELSE
      expandedKey(197);
  
  out0_111(198) <= out0_110(198) WHEN out0_20 = '0' ELSE
      expandedKey(198);
  
  out0_111(199) <= out0_110(199) WHEN out0_20 = '0' ELSE
      expandedKey(199);
  
  out0_111(200) <= out0_110(200) WHEN out0_20 = '0' ELSE
      expandedKey(200);
  
  out0_111(201) <= out0_110(201) WHEN out0_20 = '0' ELSE
      expandedKey(201);
  
  out0_111(202) <= out0_110(202) WHEN out0_20 = '0' ELSE
      expandedKey(202);
  
  out0_111(203) <= out0_110(203) WHEN out0_20 = '0' ELSE
      expandedKey(203);
  
  out0_111(204) <= out0_110(204) WHEN out0_20 = '0' ELSE
      expandedKey(204);
  
  out0_111(205) <= out0_110(205) WHEN out0_20 = '0' ELSE
      expandedKey(205);
  
  out0_111(206) <= out0_110(206) WHEN out0_20 = '0' ELSE
      expandedKey(206);
  
  out0_111(207) <= out0_110(207) WHEN out0_20 = '0' ELSE
      expandedKey(207);
  
  out0_111(208) <= out0_110(208) WHEN out0_20 = '0' ELSE
      expandedKey(208);
  
  out0_111(209) <= out0_110(209) WHEN out0_20 = '0' ELSE
      expandedKey(209);
  
  out0_111(210) <= out0_110(210) WHEN out0_20 = '0' ELSE
      expandedKey(210);
  
  out0_111(211) <= out0_110(211) WHEN out0_20 = '0' ELSE
      expandedKey(211);
  
  out0_111(212) <= out0_110(212) WHEN out0_20 = '0' ELSE
      expandedKey(212);
  
  out0_111(213) <= out0_110(213) WHEN out0_20 = '0' ELSE
      expandedKey(213);
  
  out0_111(214) <= out0_110(214) WHEN out0_20 = '0' ELSE
      expandedKey(214);
  
  out0_111(215) <= out0_110(215) WHEN out0_20 = '0' ELSE
      expandedKey(215);
  
  out0_111(216) <= out0_110(216) WHEN out0_20 = '0' ELSE
      expandedKey(216);
  
  out0_111(217) <= out0_110(217) WHEN out0_20 = '0' ELSE
      expandedKey(217);
  
  out0_111(218) <= out0_110(218) WHEN out0_20 = '0' ELSE
      expandedKey(218);
  
  out0_111(219) <= out0_110(219) WHEN out0_20 = '0' ELSE
      expandedKey(219);
  
  out0_111(220) <= out0_110(220) WHEN out0_20 = '0' ELSE
      expandedKey(220);
  
  out0_111(221) <= out0_110(221) WHEN out0_20 = '0' ELSE
      expandedKey(221);
  
  out0_111(222) <= out0_110(222) WHEN out0_20 = '0' ELSE
      expandedKey(222);
  
  out0_111(223) <= out0_110(223) WHEN out0_20 = '0' ELSE
      expandedKey(223);
  
  out0_111(224) <= out0_110(224) WHEN out0_20 = '0' ELSE
      expandedKey(224);
  
  out0_111(225) <= out0_110(225) WHEN out0_20 = '0' ELSE
      expandedKey(225);
  
  out0_111(226) <= out0_110(226) WHEN out0_20 = '0' ELSE
      expandedKey(226);
  
  out0_111(227) <= out0_110(227) WHEN out0_20 = '0' ELSE
      expandedKey(227);
  
  out0_111(228) <= out0_110(228) WHEN out0_20 = '0' ELSE
      expandedKey(228);
  
  out0_111(229) <= out0_110(229) WHEN out0_20 = '0' ELSE
      expandedKey(229);
  
  out0_111(230) <= out0_110(230) WHEN out0_20 = '0' ELSE
      expandedKey(230);
  
  out0_111(231) <= out0_110(231) WHEN out0_20 = '0' ELSE
      expandedKey(231);
  
  out0_111(232) <= out0_110(232) WHEN out0_20 = '0' ELSE
      expandedKey(232);
  
  out0_111(233) <= out0_110(233) WHEN out0_20 = '0' ELSE
      expandedKey(233);
  
  out0_111(234) <= out0_110(234) WHEN out0_20 = '0' ELSE
      expandedKey(234);
  
  out0_111(235) <= out0_110(235) WHEN out0_20 = '0' ELSE
      expandedKey(235);
  
  out0_111(236) <= out0_110(236) WHEN out0_20 = '0' ELSE
      expandedKey(236);
  
  out0_111(237) <= out0_110(237) WHEN out0_20 = '0' ELSE
      expandedKey(237);
  
  out0_111(238) <= out0_110(238) WHEN out0_20 = '0' ELSE
      expandedKey(238);
  
  out0_111(239) <= out0_110(239) WHEN out0_20 = '0' ELSE
      expandedKey(239);

  
  out0_112(0) <= out0_111(0) WHEN out0_22 = '0' ELSE
      expandedKey_5(0);
  
  out0_112(1) <= out0_111(1) WHEN out0_22 = '0' ELSE
      expandedKey_5(1);
  
  out0_112(2) <= out0_111(2) WHEN out0_22 = '0' ELSE
      expandedKey_5(2);
  
  out0_112(3) <= out0_111(3) WHEN out0_22 = '0' ELSE
      expandedKey_5(3);
  
  out0_112(4) <= out0_111(4) WHEN out0_22 = '0' ELSE
      expandedKey_5(4);
  
  out0_112(5) <= out0_111(5) WHEN out0_22 = '0' ELSE
      expandedKey_5(5);
  
  out0_112(6) <= out0_111(6) WHEN out0_22 = '0' ELSE
      expandedKey_5(6);
  
  out0_112(7) <= out0_111(7) WHEN out0_22 = '0' ELSE
      expandedKey_5(7);
  
  out0_112(8) <= out0_111(8) WHEN out0_22 = '0' ELSE
      expandedKey_5(8);
  
  out0_112(9) <= out0_111(9) WHEN out0_22 = '0' ELSE
      expandedKey_5(9);
  
  out0_112(10) <= out0_111(10) WHEN out0_22 = '0' ELSE
      expandedKey_5(10);
  
  out0_112(11) <= out0_111(11) WHEN out0_22 = '0' ELSE
      expandedKey_5(11);
  
  out0_112(12) <= out0_111(12) WHEN out0_22 = '0' ELSE
      expandedKey_5(12);
  
  out0_112(13) <= out0_111(13) WHEN out0_22 = '0' ELSE
      expandedKey_5(13);
  
  out0_112(14) <= out0_111(14) WHEN out0_22 = '0' ELSE
      expandedKey_5(14);
  
  out0_112(15) <= out0_111(15) WHEN out0_22 = '0' ELSE
      expandedKey_5(15);
  
  out0_112(16) <= out0_111(16) WHEN out0_22 = '0' ELSE
      expandedKey_5(16);
  
  out0_112(17) <= out0_111(17) WHEN out0_22 = '0' ELSE
      expandedKey_5(17);
  
  out0_112(18) <= out0_111(18) WHEN out0_22 = '0' ELSE
      expandedKey_5(18);
  
  out0_112(19) <= out0_111(19) WHEN out0_22 = '0' ELSE
      expandedKey_5(19);
  
  out0_112(20) <= out0_111(20) WHEN out0_22 = '0' ELSE
      expandedKey_5(20);
  
  out0_112(21) <= out0_111(21) WHEN out0_22 = '0' ELSE
      expandedKey_5(21);
  
  out0_112(22) <= out0_111(22) WHEN out0_22 = '0' ELSE
      expandedKey_5(22);
  
  out0_112(23) <= out0_111(23) WHEN out0_22 = '0' ELSE
      expandedKey_5(23);
  
  out0_112(24) <= out0_111(24) WHEN out0_22 = '0' ELSE
      expandedKey_5(24);
  
  out0_112(25) <= out0_111(25) WHEN out0_22 = '0' ELSE
      expandedKey_5(25);
  
  out0_112(26) <= out0_111(26) WHEN out0_22 = '0' ELSE
      expandedKey_5(26);
  
  out0_112(27) <= out0_111(27) WHEN out0_22 = '0' ELSE
      expandedKey_5(27);
  
  out0_112(28) <= out0_111(28) WHEN out0_22 = '0' ELSE
      expandedKey_5(28);
  
  out0_112(29) <= out0_111(29) WHEN out0_22 = '0' ELSE
      expandedKey_5(29);
  
  out0_112(30) <= out0_111(30) WHEN out0_22 = '0' ELSE
      expandedKey_5(30);
  
  out0_112(31) <= out0_111(31) WHEN out0_22 = '0' ELSE
      expandedKey_5(31);
  
  out0_112(32) <= out0_111(32) WHEN out0_22 = '0' ELSE
      expandedKey_5(32);
  
  out0_112(33) <= out0_111(33) WHEN out0_22 = '0' ELSE
      expandedKey_5(33);
  
  out0_112(34) <= out0_111(34) WHEN out0_22 = '0' ELSE
      expandedKey_5(34);
  
  out0_112(35) <= out0_111(35) WHEN out0_22 = '0' ELSE
      expandedKey_5(35);
  
  out0_112(36) <= out0_111(36) WHEN out0_22 = '0' ELSE
      expandedKey_5(36);
  
  out0_112(37) <= out0_111(37) WHEN out0_22 = '0' ELSE
      expandedKey_5(37);
  
  out0_112(38) <= out0_111(38) WHEN out0_22 = '0' ELSE
      expandedKey_5(38);
  
  out0_112(39) <= out0_111(39) WHEN out0_22 = '0' ELSE
      expandedKey_5(39);
  
  out0_112(40) <= out0_111(40) WHEN out0_22 = '0' ELSE
      expandedKey_5(40);
  
  out0_112(41) <= out0_111(41) WHEN out0_22 = '0' ELSE
      expandedKey_5(41);
  
  out0_112(42) <= out0_111(42) WHEN out0_22 = '0' ELSE
      expandedKey_5(42);
  
  out0_112(43) <= out0_111(43) WHEN out0_22 = '0' ELSE
      expandedKey_5(43);
  
  out0_112(44) <= out0_111(44) WHEN out0_22 = '0' ELSE
      expandedKey_5(44);
  
  out0_112(45) <= out0_111(45) WHEN out0_22 = '0' ELSE
      expandedKey_5(45);
  
  out0_112(46) <= out0_111(46) WHEN out0_22 = '0' ELSE
      expandedKey_5(46);
  
  out0_112(47) <= out0_111(47) WHEN out0_22 = '0' ELSE
      expandedKey_5(47);
  
  out0_112(48) <= out0_111(48) WHEN out0_22 = '0' ELSE
      expandedKey_5(48);
  
  out0_112(49) <= out0_111(49) WHEN out0_22 = '0' ELSE
      expandedKey_5(49);
  
  out0_112(50) <= out0_111(50) WHEN out0_22 = '0' ELSE
      expandedKey_5(50);
  
  out0_112(51) <= out0_111(51) WHEN out0_22 = '0' ELSE
      expandedKey_5(51);
  
  out0_112(52) <= out0_111(52) WHEN out0_22 = '0' ELSE
      expandedKey_5(52);
  
  out0_112(53) <= out0_111(53) WHEN out0_22 = '0' ELSE
      expandedKey_5(53);
  
  out0_112(54) <= out0_111(54) WHEN out0_22 = '0' ELSE
      expandedKey_5(54);
  
  out0_112(55) <= out0_111(55) WHEN out0_22 = '0' ELSE
      expandedKey_5(55);
  
  out0_112(56) <= out0_111(56) WHEN out0_22 = '0' ELSE
      expandedKey_5(56);
  
  out0_112(57) <= out0_111(57) WHEN out0_22 = '0' ELSE
      expandedKey_5(57);
  
  out0_112(58) <= out0_111(58) WHEN out0_22 = '0' ELSE
      expandedKey_5(58);
  
  out0_112(59) <= out0_111(59) WHEN out0_22 = '0' ELSE
      expandedKey_5(59);
  
  out0_112(60) <= out0_111(60) WHEN out0_22 = '0' ELSE
      expandedKey_5(60);
  
  out0_112(61) <= out0_111(61) WHEN out0_22 = '0' ELSE
      expandedKey_5(61);
  
  out0_112(62) <= out0_111(62) WHEN out0_22 = '0' ELSE
      expandedKey_5(62);
  
  out0_112(63) <= out0_111(63) WHEN out0_22 = '0' ELSE
      expandedKey_5(63);
  
  out0_112(64) <= out0_111(64) WHEN out0_22 = '0' ELSE
      expandedKey_5(64);
  
  out0_112(65) <= out0_111(65) WHEN out0_22 = '0' ELSE
      expandedKey_5(65);
  
  out0_112(66) <= out0_111(66) WHEN out0_22 = '0' ELSE
      expandedKey_5(66);
  
  out0_112(67) <= out0_111(67) WHEN out0_22 = '0' ELSE
      expandedKey_5(67);
  
  out0_112(68) <= out0_111(68) WHEN out0_22 = '0' ELSE
      expandedKey_5(68);
  
  out0_112(69) <= out0_111(69) WHEN out0_22 = '0' ELSE
      expandedKey_5(69);
  
  out0_112(70) <= out0_111(70) WHEN out0_22 = '0' ELSE
      expandedKey_5(70);
  
  out0_112(71) <= out0_111(71) WHEN out0_22 = '0' ELSE
      expandedKey_5(71);
  
  out0_112(72) <= out0_111(72) WHEN out0_22 = '0' ELSE
      expandedKey_5(72);
  
  out0_112(73) <= out0_111(73) WHEN out0_22 = '0' ELSE
      expandedKey_5(73);
  
  out0_112(74) <= out0_111(74) WHEN out0_22 = '0' ELSE
      expandedKey_5(74);
  
  out0_112(75) <= out0_111(75) WHEN out0_22 = '0' ELSE
      expandedKey_5(75);
  
  out0_112(76) <= out0_111(76) WHEN out0_22 = '0' ELSE
      expandedKey_5(76);
  
  out0_112(77) <= out0_111(77) WHEN out0_22 = '0' ELSE
      expandedKey_5(77);
  
  out0_112(78) <= out0_111(78) WHEN out0_22 = '0' ELSE
      expandedKey_5(78);
  
  out0_112(79) <= out0_111(79) WHEN out0_22 = '0' ELSE
      expandedKey_5(79);
  
  out0_112(80) <= out0_111(80) WHEN out0_22 = '0' ELSE
      expandedKey_5(80);
  
  out0_112(81) <= out0_111(81) WHEN out0_22 = '0' ELSE
      expandedKey_5(81);
  
  out0_112(82) <= out0_111(82) WHEN out0_22 = '0' ELSE
      expandedKey_5(82);
  
  out0_112(83) <= out0_111(83) WHEN out0_22 = '0' ELSE
      expandedKey_5(83);
  
  out0_112(84) <= out0_111(84) WHEN out0_22 = '0' ELSE
      expandedKey_5(84);
  
  out0_112(85) <= out0_111(85) WHEN out0_22 = '0' ELSE
      expandedKey_5(85);
  
  out0_112(86) <= out0_111(86) WHEN out0_22 = '0' ELSE
      expandedKey_5(86);
  
  out0_112(87) <= out0_111(87) WHEN out0_22 = '0' ELSE
      expandedKey_5(87);
  
  out0_112(88) <= out0_111(88) WHEN out0_22 = '0' ELSE
      expandedKey_5(88);
  
  out0_112(89) <= out0_111(89) WHEN out0_22 = '0' ELSE
      expandedKey_5(89);
  
  out0_112(90) <= out0_111(90) WHEN out0_22 = '0' ELSE
      expandedKey_5(90);
  
  out0_112(91) <= out0_111(91) WHEN out0_22 = '0' ELSE
      expandedKey_5(91);
  
  out0_112(92) <= out0_111(92) WHEN out0_22 = '0' ELSE
      expandedKey_5(92);
  
  out0_112(93) <= out0_111(93) WHEN out0_22 = '0' ELSE
      expandedKey_5(93);
  
  out0_112(94) <= out0_111(94) WHEN out0_22 = '0' ELSE
      expandedKey_5(94);
  
  out0_112(95) <= out0_111(95) WHEN out0_22 = '0' ELSE
      expandedKey_5(95);
  
  out0_112(96) <= out0_111(96) WHEN out0_22 = '0' ELSE
      expandedKey_5(96);
  
  out0_112(97) <= out0_111(97) WHEN out0_22 = '0' ELSE
      expandedKey_5(97);
  
  out0_112(98) <= out0_111(98) WHEN out0_22 = '0' ELSE
      expandedKey_5(98);
  
  out0_112(99) <= out0_111(99) WHEN out0_22 = '0' ELSE
      expandedKey_5(99);
  
  out0_112(100) <= out0_111(100) WHEN out0_22 = '0' ELSE
      expandedKey_5(100);
  
  out0_112(101) <= out0_111(101) WHEN out0_22 = '0' ELSE
      expandedKey_5(101);
  
  out0_112(102) <= out0_111(102) WHEN out0_22 = '0' ELSE
      expandedKey_5(102);
  
  out0_112(103) <= out0_111(103) WHEN out0_22 = '0' ELSE
      expandedKey_5(103);
  
  out0_112(104) <= out0_111(104) WHEN out0_22 = '0' ELSE
      expandedKey_5(104);
  
  out0_112(105) <= out0_111(105) WHEN out0_22 = '0' ELSE
      expandedKey_5(105);
  
  out0_112(106) <= out0_111(106) WHEN out0_22 = '0' ELSE
      expandedKey_5(106);
  
  out0_112(107) <= out0_111(107) WHEN out0_22 = '0' ELSE
      expandedKey_5(107);
  
  out0_112(108) <= out0_111(108) WHEN out0_22 = '0' ELSE
      expandedKey_5(108);
  
  out0_112(109) <= out0_111(109) WHEN out0_22 = '0' ELSE
      expandedKey_5(109);
  
  out0_112(110) <= out0_111(110) WHEN out0_22 = '0' ELSE
      expandedKey_5(110);
  
  out0_112(111) <= out0_111(111) WHEN out0_22 = '0' ELSE
      expandedKey_5(111);
  
  out0_112(112) <= out0_111(112) WHEN out0_22 = '0' ELSE
      expandedKey_5(112);
  
  out0_112(113) <= out0_111(113) WHEN out0_22 = '0' ELSE
      expandedKey_5(113);
  
  out0_112(114) <= out0_111(114) WHEN out0_22 = '0' ELSE
      expandedKey_5(114);
  
  out0_112(115) <= out0_111(115) WHEN out0_22 = '0' ELSE
      expandedKey_5(115);
  
  out0_112(116) <= out0_111(116) WHEN out0_22 = '0' ELSE
      expandedKey_5(116);
  
  out0_112(117) <= out0_111(117) WHEN out0_22 = '0' ELSE
      expandedKey_5(117);
  
  out0_112(118) <= out0_111(118) WHEN out0_22 = '0' ELSE
      expandedKey_5(118);
  
  out0_112(119) <= out0_111(119) WHEN out0_22 = '0' ELSE
      expandedKey_5(119);
  
  out0_112(120) <= out0_111(120) WHEN out0_22 = '0' ELSE
      expandedKey_5(120);
  
  out0_112(121) <= out0_111(121) WHEN out0_22 = '0' ELSE
      expandedKey_5(121);
  
  out0_112(122) <= out0_111(122) WHEN out0_22 = '0' ELSE
      expandedKey_5(122);
  
  out0_112(123) <= out0_111(123) WHEN out0_22 = '0' ELSE
      expandedKey_5(123);
  
  out0_112(124) <= out0_111(124) WHEN out0_22 = '0' ELSE
      expandedKey_5(124);
  
  out0_112(125) <= out0_111(125) WHEN out0_22 = '0' ELSE
      expandedKey_5(125);
  
  out0_112(126) <= out0_111(126) WHEN out0_22 = '0' ELSE
      expandedKey_5(126);
  
  out0_112(127) <= out0_111(127) WHEN out0_22 = '0' ELSE
      expandedKey_5(127);
  
  out0_112(128) <= out0_111(128) WHEN out0_22 = '0' ELSE
      expandedKey_5(128);
  
  out0_112(129) <= out0_111(129) WHEN out0_22 = '0' ELSE
      expandedKey_5(129);
  
  out0_112(130) <= out0_111(130) WHEN out0_22 = '0' ELSE
      expandedKey_5(130);
  
  out0_112(131) <= out0_111(131) WHEN out0_22 = '0' ELSE
      expandedKey_5(131);
  
  out0_112(132) <= out0_111(132) WHEN out0_22 = '0' ELSE
      expandedKey_5(132);
  
  out0_112(133) <= out0_111(133) WHEN out0_22 = '0' ELSE
      expandedKey_5(133);
  
  out0_112(134) <= out0_111(134) WHEN out0_22 = '0' ELSE
      expandedKey_5(134);
  
  out0_112(135) <= out0_111(135) WHEN out0_22 = '0' ELSE
      expandedKey_5(135);
  
  out0_112(136) <= out0_111(136) WHEN out0_22 = '0' ELSE
      expandedKey_5(136);
  
  out0_112(137) <= out0_111(137) WHEN out0_22 = '0' ELSE
      expandedKey_5(137);
  
  out0_112(138) <= out0_111(138) WHEN out0_22 = '0' ELSE
      expandedKey_5(138);
  
  out0_112(139) <= out0_111(139) WHEN out0_22 = '0' ELSE
      expandedKey_5(139);
  
  out0_112(140) <= out0_111(140) WHEN out0_22 = '0' ELSE
      expandedKey_5(140);
  
  out0_112(141) <= out0_111(141) WHEN out0_22 = '0' ELSE
      expandedKey_5(141);
  
  out0_112(142) <= out0_111(142) WHEN out0_22 = '0' ELSE
      expandedKey_5(142);
  
  out0_112(143) <= out0_111(143) WHEN out0_22 = '0' ELSE
      expandedKey_5(143);
  
  out0_112(144) <= out0_111(144) WHEN out0_22 = '0' ELSE
      expandedKey_5(144);
  
  out0_112(145) <= out0_111(145) WHEN out0_22 = '0' ELSE
      expandedKey_5(145);
  
  out0_112(146) <= out0_111(146) WHEN out0_22 = '0' ELSE
      expandedKey_5(146);
  
  out0_112(147) <= out0_111(147) WHEN out0_22 = '0' ELSE
      expandedKey_5(147);
  
  out0_112(148) <= out0_111(148) WHEN out0_22 = '0' ELSE
      expandedKey_5(148);
  
  out0_112(149) <= out0_111(149) WHEN out0_22 = '0' ELSE
      expandedKey_5(149);
  
  out0_112(150) <= out0_111(150) WHEN out0_22 = '0' ELSE
      expandedKey_5(150);
  
  out0_112(151) <= out0_111(151) WHEN out0_22 = '0' ELSE
      expandedKey_5(151);
  
  out0_112(152) <= out0_111(152) WHEN out0_22 = '0' ELSE
      expandedKey_5(152);
  
  out0_112(153) <= out0_111(153) WHEN out0_22 = '0' ELSE
      expandedKey_5(153);
  
  out0_112(154) <= out0_111(154) WHEN out0_22 = '0' ELSE
      expandedKey_5(154);
  
  out0_112(155) <= out0_111(155) WHEN out0_22 = '0' ELSE
      expandedKey_5(155);
  
  out0_112(156) <= out0_111(156) WHEN out0_22 = '0' ELSE
      expandedKey_5(156);
  
  out0_112(157) <= out0_111(157) WHEN out0_22 = '0' ELSE
      expandedKey_5(157);
  
  out0_112(158) <= out0_111(158) WHEN out0_22 = '0' ELSE
      expandedKey_5(158);
  
  out0_112(159) <= out0_111(159) WHEN out0_22 = '0' ELSE
      expandedKey_5(159);
  
  out0_112(160) <= out0_111(160) WHEN out0_22 = '0' ELSE
      expandedKey_5(160);
  
  out0_112(161) <= out0_111(161) WHEN out0_22 = '0' ELSE
      expandedKey_5(161);
  
  out0_112(162) <= out0_111(162) WHEN out0_22 = '0' ELSE
      expandedKey_5(162);
  
  out0_112(163) <= out0_111(163) WHEN out0_22 = '0' ELSE
      expandedKey_5(163);
  
  out0_112(164) <= out0_111(164) WHEN out0_22 = '0' ELSE
      expandedKey_5(164);
  
  out0_112(165) <= out0_111(165) WHEN out0_22 = '0' ELSE
      expandedKey_5(165);
  
  out0_112(166) <= out0_111(166) WHEN out0_22 = '0' ELSE
      expandedKey_5(166);
  
  out0_112(167) <= out0_111(167) WHEN out0_22 = '0' ELSE
      expandedKey_5(167);
  
  out0_112(168) <= out0_111(168) WHEN out0_22 = '0' ELSE
      expandedKey_5(168);
  
  out0_112(169) <= out0_111(169) WHEN out0_22 = '0' ELSE
      expandedKey_5(169);
  
  out0_112(170) <= out0_111(170) WHEN out0_22 = '0' ELSE
      expandedKey_5(170);
  
  out0_112(171) <= out0_111(171) WHEN out0_22 = '0' ELSE
      expandedKey_5(171);
  
  out0_112(172) <= out0_111(172) WHEN out0_22 = '0' ELSE
      expandedKey_5(172);
  
  out0_112(173) <= out0_111(173) WHEN out0_22 = '0' ELSE
      expandedKey_5(173);
  
  out0_112(174) <= out0_111(174) WHEN out0_22 = '0' ELSE
      expandedKey_5(174);
  
  out0_112(175) <= out0_111(175) WHEN out0_22 = '0' ELSE
      expandedKey_5(175);
  
  out0_112(176) <= out0_111(176) WHEN out0_22 = '0' ELSE
      expandedKey_5(176);
  
  out0_112(177) <= out0_111(177) WHEN out0_22 = '0' ELSE
      expandedKey_5(177);
  
  out0_112(178) <= out0_111(178) WHEN out0_22 = '0' ELSE
      expandedKey_5(178);
  
  out0_112(179) <= out0_111(179) WHEN out0_22 = '0' ELSE
      expandedKey_5(179);
  
  out0_112(180) <= out0_111(180) WHEN out0_22 = '0' ELSE
      expandedKey_5(180);
  
  out0_112(181) <= out0_111(181) WHEN out0_22 = '0' ELSE
      expandedKey_5(181);
  
  out0_112(182) <= out0_111(182) WHEN out0_22 = '0' ELSE
      expandedKey_5(182);
  
  out0_112(183) <= out0_111(183) WHEN out0_22 = '0' ELSE
      expandedKey_5(183);
  
  out0_112(184) <= out0_111(184) WHEN out0_22 = '0' ELSE
      expandedKey_5(184);
  
  out0_112(185) <= out0_111(185) WHEN out0_22 = '0' ELSE
      expandedKey_5(185);
  
  out0_112(186) <= out0_111(186) WHEN out0_22 = '0' ELSE
      expandedKey_5(186);
  
  out0_112(187) <= out0_111(187) WHEN out0_22 = '0' ELSE
      expandedKey_5(187);
  
  out0_112(188) <= out0_111(188) WHEN out0_22 = '0' ELSE
      expandedKey_5(188);
  
  out0_112(189) <= out0_111(189) WHEN out0_22 = '0' ELSE
      expandedKey_5(189);
  
  out0_112(190) <= out0_111(190) WHEN out0_22 = '0' ELSE
      expandedKey_5(190);
  
  out0_112(191) <= out0_111(191) WHEN out0_22 = '0' ELSE
      expandedKey_5(191);
  
  out0_112(192) <= out0_111(192) WHEN out0_22 = '0' ELSE
      expandedKey_5(192);
  
  out0_112(193) <= out0_111(193) WHEN out0_22 = '0' ELSE
      expandedKey_5(193);
  
  out0_112(194) <= out0_111(194) WHEN out0_22 = '0' ELSE
      expandedKey_5(194);
  
  out0_112(195) <= out0_111(195) WHEN out0_22 = '0' ELSE
      expandedKey_5(195);
  
  out0_112(196) <= out0_111(196) WHEN out0_22 = '0' ELSE
      expandedKey_5(196);
  
  out0_112(197) <= out0_111(197) WHEN out0_22 = '0' ELSE
      expandedKey_5(197);
  
  out0_112(198) <= out0_111(198) WHEN out0_22 = '0' ELSE
      expandedKey_5(198);
  
  out0_112(199) <= out0_111(199) WHEN out0_22 = '0' ELSE
      expandedKey_5(199);
  
  out0_112(200) <= out0_111(200) WHEN out0_22 = '0' ELSE
      expandedKey_5(200);
  
  out0_112(201) <= out0_111(201) WHEN out0_22 = '0' ELSE
      expandedKey_5(201);
  
  out0_112(202) <= out0_111(202) WHEN out0_22 = '0' ELSE
      expandedKey_5(202);
  
  out0_112(203) <= out0_111(203) WHEN out0_22 = '0' ELSE
      expandedKey_5(203);
  
  out0_112(204) <= out0_111(204) WHEN out0_22 = '0' ELSE
      expandedKey_5(204);
  
  out0_112(205) <= out0_111(205) WHEN out0_22 = '0' ELSE
      expandedKey_5(205);
  
  out0_112(206) <= out0_111(206) WHEN out0_22 = '0' ELSE
      expandedKey_5(206);
  
  out0_112(207) <= out0_111(207) WHEN out0_22 = '0' ELSE
      expandedKey_5(207);
  
  out0_112(208) <= out0_111(208) WHEN out0_22 = '0' ELSE
      expandedKey_5(208);
  
  out0_112(209) <= out0_111(209) WHEN out0_22 = '0' ELSE
      expandedKey_5(209);
  
  out0_112(210) <= out0_111(210) WHEN out0_22 = '0' ELSE
      expandedKey_5(210);
  
  out0_112(211) <= out0_111(211) WHEN out0_22 = '0' ELSE
      expandedKey_5(211);
  
  out0_112(212) <= out0_111(212) WHEN out0_22 = '0' ELSE
      expandedKey_5(212);
  
  out0_112(213) <= out0_111(213) WHEN out0_22 = '0' ELSE
      expandedKey_5(213);
  
  out0_112(214) <= out0_111(214) WHEN out0_22 = '0' ELSE
      expandedKey_5(214);
  
  out0_112(215) <= out0_111(215) WHEN out0_22 = '0' ELSE
      expandedKey_5(215);
  
  out0_112(216) <= out0_111(216) WHEN out0_22 = '0' ELSE
      expandedKey_5(216);
  
  out0_112(217) <= out0_111(217) WHEN out0_22 = '0' ELSE
      expandedKey_5(217);
  
  out0_112(218) <= out0_111(218) WHEN out0_22 = '0' ELSE
      expandedKey_5(218);
  
  out0_112(219) <= out0_111(219) WHEN out0_22 = '0' ELSE
      expandedKey_5(219);
  
  out0_112(220) <= out0_111(220) WHEN out0_22 = '0' ELSE
      expandedKey_5(220);
  
  out0_112(221) <= out0_111(221) WHEN out0_22 = '0' ELSE
      expandedKey_5(221);
  
  out0_112(222) <= out0_111(222) WHEN out0_22 = '0' ELSE
      expandedKey_5(222);
  
  out0_112(223) <= out0_111(223) WHEN out0_22 = '0' ELSE
      expandedKey_5(223);
  
  out0_112(224) <= out0_111(224) WHEN out0_22 = '0' ELSE
      expandedKey_5(224);
  
  out0_112(225) <= out0_111(225) WHEN out0_22 = '0' ELSE
      expandedKey_5(225);
  
  out0_112(226) <= out0_111(226) WHEN out0_22 = '0' ELSE
      expandedKey_5(226);
  
  out0_112(227) <= out0_111(227) WHEN out0_22 = '0' ELSE
      expandedKey_5(227);
  
  out0_112(228) <= out0_111(228) WHEN out0_22 = '0' ELSE
      expandedKey_5(228);
  
  out0_112(229) <= out0_111(229) WHEN out0_22 = '0' ELSE
      expandedKey_5(229);
  
  out0_112(230) <= out0_111(230) WHEN out0_22 = '0' ELSE
      expandedKey_5(230);
  
  out0_112(231) <= out0_111(231) WHEN out0_22 = '0' ELSE
      expandedKey_5(231);
  
  out0_112(232) <= out0_111(232) WHEN out0_22 = '0' ELSE
      expandedKey_5(232);
  
  out0_112(233) <= out0_111(233) WHEN out0_22 = '0' ELSE
      expandedKey_5(233);
  
  out0_112(234) <= out0_111(234) WHEN out0_22 = '0' ELSE
      expandedKey_5(234);
  
  out0_112(235) <= out0_111(235) WHEN out0_22 = '0' ELSE
      expandedKey_5(235);
  
  out0_112(236) <= out0_111(236) WHEN out0_22 = '0' ELSE
      expandedKey_5(236);
  
  out0_112(237) <= out0_111(237) WHEN out0_22 = '0' ELSE
      expandedKey_5(237);
  
  out0_112(238) <= out0_111(238) WHEN out0_22 = '0' ELSE
      expandedKey_5(238);
  
  out0_112(239) <= out0_111(239) WHEN out0_22 = '0' ELSE
      expandedKey_5(239);

  
  expandedKey_6(0) <= out0_112(0) WHEN out0_24 = '0' ELSE
      expandedKey_1(0);
  
  expandedKey_6(1) <= out0_112(1) WHEN out0_24 = '0' ELSE
      expandedKey_1(1);
  
  expandedKey_6(2) <= out0_112(2) WHEN out0_24 = '0' ELSE
      expandedKey_1(2);
  
  expandedKey_6(3) <= out0_112(3) WHEN out0_24 = '0' ELSE
      expandedKey_1(3);
  
  expandedKey_6(4) <= out0_112(4) WHEN out0_24 = '0' ELSE
      expandedKey_1(4);
  
  expandedKey_6(5) <= out0_112(5) WHEN out0_24 = '0' ELSE
      expandedKey_1(5);
  
  expandedKey_6(6) <= out0_112(6) WHEN out0_24 = '0' ELSE
      expandedKey_1(6);
  
  expandedKey_6(7) <= out0_112(7) WHEN out0_24 = '0' ELSE
      expandedKey_1(7);
  
  expandedKey_6(8) <= out0_112(8) WHEN out0_24 = '0' ELSE
      expandedKey_1(8);
  
  expandedKey_6(9) <= out0_112(9) WHEN out0_24 = '0' ELSE
      expandedKey_1(9);
  
  expandedKey_6(10) <= out0_112(10) WHEN out0_24 = '0' ELSE
      expandedKey_1(10);
  
  expandedKey_6(11) <= out0_112(11) WHEN out0_24 = '0' ELSE
      expandedKey_1(11);
  
  expandedKey_6(12) <= out0_112(12) WHEN out0_24 = '0' ELSE
      expandedKey_1(12);
  
  expandedKey_6(13) <= out0_112(13) WHEN out0_24 = '0' ELSE
      expandedKey_1(13);
  
  expandedKey_6(14) <= out0_112(14) WHEN out0_24 = '0' ELSE
      expandedKey_1(14);
  
  expandedKey_6(15) <= out0_112(15) WHEN out0_24 = '0' ELSE
      expandedKey_1(15);
  
  expandedKey_6(16) <= out0_112(16) WHEN out0_24 = '0' ELSE
      expandedKey_1(16);
  
  expandedKey_6(17) <= out0_112(17) WHEN out0_24 = '0' ELSE
      expandedKey_1(17);
  
  expandedKey_6(18) <= out0_112(18) WHEN out0_24 = '0' ELSE
      expandedKey_1(18);
  
  expandedKey_6(19) <= out0_112(19) WHEN out0_24 = '0' ELSE
      expandedKey_1(19);
  
  expandedKey_6(20) <= out0_112(20) WHEN out0_24 = '0' ELSE
      expandedKey_1(20);
  
  expandedKey_6(21) <= out0_112(21) WHEN out0_24 = '0' ELSE
      expandedKey_1(21);
  
  expandedKey_6(22) <= out0_112(22) WHEN out0_24 = '0' ELSE
      expandedKey_1(22);
  
  expandedKey_6(23) <= out0_112(23) WHEN out0_24 = '0' ELSE
      expandedKey_1(23);
  
  expandedKey_6(24) <= out0_112(24) WHEN out0_24 = '0' ELSE
      expandedKey_1(24);
  
  expandedKey_6(25) <= out0_112(25) WHEN out0_24 = '0' ELSE
      expandedKey_1(25);
  
  expandedKey_6(26) <= out0_112(26) WHEN out0_24 = '0' ELSE
      expandedKey_1(26);
  
  expandedKey_6(27) <= out0_112(27) WHEN out0_24 = '0' ELSE
      expandedKey_1(27);
  
  expandedKey_6(28) <= out0_112(28) WHEN out0_24 = '0' ELSE
      expandedKey_1(28);
  
  expandedKey_6(29) <= out0_112(29) WHEN out0_24 = '0' ELSE
      expandedKey_1(29);
  
  expandedKey_6(30) <= out0_112(30) WHEN out0_24 = '0' ELSE
      expandedKey_1(30);
  
  expandedKey_6(31) <= out0_112(31) WHEN out0_24 = '0' ELSE
      expandedKey_1(31);
  
  expandedKey_6(32) <= out0_112(32) WHEN out0_24 = '0' ELSE
      expandedKey_1(32);
  
  expandedKey_6(33) <= out0_112(33) WHEN out0_24 = '0' ELSE
      expandedKey_1(33);
  
  expandedKey_6(34) <= out0_112(34) WHEN out0_24 = '0' ELSE
      expandedKey_1(34);
  
  expandedKey_6(35) <= out0_112(35) WHEN out0_24 = '0' ELSE
      expandedKey_1(35);
  
  expandedKey_6(36) <= out0_112(36) WHEN out0_24 = '0' ELSE
      expandedKey_1(36);
  
  expandedKey_6(37) <= out0_112(37) WHEN out0_24 = '0' ELSE
      expandedKey_1(37);
  
  expandedKey_6(38) <= out0_112(38) WHEN out0_24 = '0' ELSE
      expandedKey_1(38);
  
  expandedKey_6(39) <= out0_112(39) WHEN out0_24 = '0' ELSE
      expandedKey_1(39);
  
  expandedKey_6(40) <= out0_112(40) WHEN out0_24 = '0' ELSE
      expandedKey_1(40);
  
  expandedKey_6(41) <= out0_112(41) WHEN out0_24 = '0' ELSE
      expandedKey_1(41);
  
  expandedKey_6(42) <= out0_112(42) WHEN out0_24 = '0' ELSE
      expandedKey_1(42);
  
  expandedKey_6(43) <= out0_112(43) WHEN out0_24 = '0' ELSE
      expandedKey_1(43);
  
  expandedKey_6(44) <= out0_112(44) WHEN out0_24 = '0' ELSE
      expandedKey_1(44);
  
  expandedKey_6(45) <= out0_112(45) WHEN out0_24 = '0' ELSE
      expandedKey_1(45);
  
  expandedKey_6(46) <= out0_112(46) WHEN out0_24 = '0' ELSE
      expandedKey_1(46);
  
  expandedKey_6(47) <= out0_112(47) WHEN out0_24 = '0' ELSE
      expandedKey_1(47);
  
  expandedKey_6(48) <= out0_112(48) WHEN out0_24 = '0' ELSE
      expandedKey_1(48);
  
  expandedKey_6(49) <= out0_112(49) WHEN out0_24 = '0' ELSE
      expandedKey_1(49);
  
  expandedKey_6(50) <= out0_112(50) WHEN out0_24 = '0' ELSE
      expandedKey_1(50);
  
  expandedKey_6(51) <= out0_112(51) WHEN out0_24 = '0' ELSE
      expandedKey_1(51);
  
  expandedKey_6(52) <= out0_112(52) WHEN out0_24 = '0' ELSE
      expandedKey_1(52);
  
  expandedKey_6(53) <= out0_112(53) WHEN out0_24 = '0' ELSE
      expandedKey_1(53);
  
  expandedKey_6(54) <= out0_112(54) WHEN out0_24 = '0' ELSE
      expandedKey_1(54);
  
  expandedKey_6(55) <= out0_112(55) WHEN out0_24 = '0' ELSE
      expandedKey_1(55);
  
  expandedKey_6(56) <= out0_112(56) WHEN out0_24 = '0' ELSE
      expandedKey_1(56);
  
  expandedKey_6(57) <= out0_112(57) WHEN out0_24 = '0' ELSE
      expandedKey_1(57);
  
  expandedKey_6(58) <= out0_112(58) WHEN out0_24 = '0' ELSE
      expandedKey_1(58);
  
  expandedKey_6(59) <= out0_112(59) WHEN out0_24 = '0' ELSE
      expandedKey_1(59);
  
  expandedKey_6(60) <= out0_112(60) WHEN out0_24 = '0' ELSE
      expandedKey_1(60);
  
  expandedKey_6(61) <= out0_112(61) WHEN out0_24 = '0' ELSE
      expandedKey_1(61);
  
  expandedKey_6(62) <= out0_112(62) WHEN out0_24 = '0' ELSE
      expandedKey_1(62);
  
  expandedKey_6(63) <= out0_112(63) WHEN out0_24 = '0' ELSE
      expandedKey_1(63);
  
  expandedKey_6(64) <= out0_112(64) WHEN out0_24 = '0' ELSE
      expandedKey_1(64);
  
  expandedKey_6(65) <= out0_112(65) WHEN out0_24 = '0' ELSE
      expandedKey_1(65);
  
  expandedKey_6(66) <= out0_112(66) WHEN out0_24 = '0' ELSE
      expandedKey_1(66);
  
  expandedKey_6(67) <= out0_112(67) WHEN out0_24 = '0' ELSE
      expandedKey_1(67);
  
  expandedKey_6(68) <= out0_112(68) WHEN out0_24 = '0' ELSE
      expandedKey_1(68);
  
  expandedKey_6(69) <= out0_112(69) WHEN out0_24 = '0' ELSE
      expandedKey_1(69);
  
  expandedKey_6(70) <= out0_112(70) WHEN out0_24 = '0' ELSE
      expandedKey_1(70);
  
  expandedKey_6(71) <= out0_112(71) WHEN out0_24 = '0' ELSE
      expandedKey_1(71);
  
  expandedKey_6(72) <= out0_112(72) WHEN out0_24 = '0' ELSE
      expandedKey_1(72);
  
  expandedKey_6(73) <= out0_112(73) WHEN out0_24 = '0' ELSE
      expandedKey_1(73);
  
  expandedKey_6(74) <= out0_112(74) WHEN out0_24 = '0' ELSE
      expandedKey_1(74);
  
  expandedKey_6(75) <= out0_112(75) WHEN out0_24 = '0' ELSE
      expandedKey_1(75);
  
  expandedKey_6(76) <= out0_112(76) WHEN out0_24 = '0' ELSE
      expandedKey_1(76);
  
  expandedKey_6(77) <= out0_112(77) WHEN out0_24 = '0' ELSE
      expandedKey_1(77);
  
  expandedKey_6(78) <= out0_112(78) WHEN out0_24 = '0' ELSE
      expandedKey_1(78);
  
  expandedKey_6(79) <= out0_112(79) WHEN out0_24 = '0' ELSE
      expandedKey_1(79);
  
  expandedKey_6(80) <= out0_112(80) WHEN out0_24 = '0' ELSE
      expandedKey_1(80);
  
  expandedKey_6(81) <= out0_112(81) WHEN out0_24 = '0' ELSE
      expandedKey_1(81);
  
  expandedKey_6(82) <= out0_112(82) WHEN out0_24 = '0' ELSE
      expandedKey_1(82);
  
  expandedKey_6(83) <= out0_112(83) WHEN out0_24 = '0' ELSE
      expandedKey_1(83);
  
  expandedKey_6(84) <= out0_112(84) WHEN out0_24 = '0' ELSE
      expandedKey_1(84);
  
  expandedKey_6(85) <= out0_112(85) WHEN out0_24 = '0' ELSE
      expandedKey_1(85);
  
  expandedKey_6(86) <= out0_112(86) WHEN out0_24 = '0' ELSE
      expandedKey_1(86);
  
  expandedKey_6(87) <= out0_112(87) WHEN out0_24 = '0' ELSE
      expandedKey_1(87);
  
  expandedKey_6(88) <= out0_112(88) WHEN out0_24 = '0' ELSE
      expandedKey_1(88);
  
  expandedKey_6(89) <= out0_112(89) WHEN out0_24 = '0' ELSE
      expandedKey_1(89);
  
  expandedKey_6(90) <= out0_112(90) WHEN out0_24 = '0' ELSE
      expandedKey_1(90);
  
  expandedKey_6(91) <= out0_112(91) WHEN out0_24 = '0' ELSE
      expandedKey_1(91);
  
  expandedKey_6(92) <= out0_112(92) WHEN out0_24 = '0' ELSE
      expandedKey_1(92);
  
  expandedKey_6(93) <= out0_112(93) WHEN out0_24 = '0' ELSE
      expandedKey_1(93);
  
  expandedKey_6(94) <= out0_112(94) WHEN out0_24 = '0' ELSE
      expandedKey_1(94);
  
  expandedKey_6(95) <= out0_112(95) WHEN out0_24 = '0' ELSE
      expandedKey_1(95);
  
  expandedKey_6(96) <= out0_112(96) WHEN out0_24 = '0' ELSE
      expandedKey_1(96);
  
  expandedKey_6(97) <= out0_112(97) WHEN out0_24 = '0' ELSE
      expandedKey_1(97);
  
  expandedKey_6(98) <= out0_112(98) WHEN out0_24 = '0' ELSE
      expandedKey_1(98);
  
  expandedKey_6(99) <= out0_112(99) WHEN out0_24 = '0' ELSE
      expandedKey_1(99);
  
  expandedKey_6(100) <= out0_112(100) WHEN out0_24 = '0' ELSE
      expandedKey_1(100);
  
  expandedKey_6(101) <= out0_112(101) WHEN out0_24 = '0' ELSE
      expandedKey_1(101);
  
  expandedKey_6(102) <= out0_112(102) WHEN out0_24 = '0' ELSE
      expandedKey_1(102);
  
  expandedKey_6(103) <= out0_112(103) WHEN out0_24 = '0' ELSE
      expandedKey_1(103);
  
  expandedKey_6(104) <= out0_112(104) WHEN out0_24 = '0' ELSE
      expandedKey_1(104);
  
  expandedKey_6(105) <= out0_112(105) WHEN out0_24 = '0' ELSE
      expandedKey_1(105);
  
  expandedKey_6(106) <= out0_112(106) WHEN out0_24 = '0' ELSE
      expandedKey_1(106);
  
  expandedKey_6(107) <= out0_112(107) WHEN out0_24 = '0' ELSE
      expandedKey_1(107);
  
  expandedKey_6(108) <= out0_112(108) WHEN out0_24 = '0' ELSE
      expandedKey_1(108);
  
  expandedKey_6(109) <= out0_112(109) WHEN out0_24 = '0' ELSE
      expandedKey_1(109);
  
  expandedKey_6(110) <= out0_112(110) WHEN out0_24 = '0' ELSE
      expandedKey_1(110);
  
  expandedKey_6(111) <= out0_112(111) WHEN out0_24 = '0' ELSE
      expandedKey_1(111);
  
  expandedKey_6(112) <= out0_112(112) WHEN out0_24 = '0' ELSE
      expandedKey_1(112);
  
  expandedKey_6(113) <= out0_112(113) WHEN out0_24 = '0' ELSE
      expandedKey_1(113);
  
  expandedKey_6(114) <= out0_112(114) WHEN out0_24 = '0' ELSE
      expandedKey_1(114);
  
  expandedKey_6(115) <= out0_112(115) WHEN out0_24 = '0' ELSE
      expandedKey_1(115);
  
  expandedKey_6(116) <= out0_112(116) WHEN out0_24 = '0' ELSE
      expandedKey_1(116);
  
  expandedKey_6(117) <= out0_112(117) WHEN out0_24 = '0' ELSE
      expandedKey_1(117);
  
  expandedKey_6(118) <= out0_112(118) WHEN out0_24 = '0' ELSE
      expandedKey_1(118);
  
  expandedKey_6(119) <= out0_112(119) WHEN out0_24 = '0' ELSE
      expandedKey_1(119);
  
  expandedKey_6(120) <= out0_112(120) WHEN out0_24 = '0' ELSE
      expandedKey_1(120);
  
  expandedKey_6(121) <= out0_112(121) WHEN out0_24 = '0' ELSE
      expandedKey_1(121);
  
  expandedKey_6(122) <= out0_112(122) WHEN out0_24 = '0' ELSE
      expandedKey_1(122);
  
  expandedKey_6(123) <= out0_112(123) WHEN out0_24 = '0' ELSE
      expandedKey_1(123);
  
  expandedKey_6(124) <= out0_112(124) WHEN out0_24 = '0' ELSE
      expandedKey_1(124);
  
  expandedKey_6(125) <= out0_112(125) WHEN out0_24 = '0' ELSE
      expandedKey_1(125);
  
  expandedKey_6(126) <= out0_112(126) WHEN out0_24 = '0' ELSE
      expandedKey_1(126);
  
  expandedKey_6(127) <= out0_112(127) WHEN out0_24 = '0' ELSE
      expandedKey_1(127);
  
  expandedKey_6(128) <= out0_112(128) WHEN out0_24 = '0' ELSE
      expandedKey_1(128);
  
  expandedKey_6(129) <= out0_112(129) WHEN out0_24 = '0' ELSE
      expandedKey_1(129);
  
  expandedKey_6(130) <= out0_112(130) WHEN out0_24 = '0' ELSE
      expandedKey_1(130);
  
  expandedKey_6(131) <= out0_112(131) WHEN out0_24 = '0' ELSE
      expandedKey_1(131);
  
  expandedKey_6(132) <= out0_112(132) WHEN out0_24 = '0' ELSE
      expandedKey_1(132);
  
  expandedKey_6(133) <= out0_112(133) WHEN out0_24 = '0' ELSE
      expandedKey_1(133);
  
  expandedKey_6(134) <= out0_112(134) WHEN out0_24 = '0' ELSE
      expandedKey_1(134);
  
  expandedKey_6(135) <= out0_112(135) WHEN out0_24 = '0' ELSE
      expandedKey_1(135);
  
  expandedKey_6(136) <= out0_112(136) WHEN out0_24 = '0' ELSE
      expandedKey_1(136);
  
  expandedKey_6(137) <= out0_112(137) WHEN out0_24 = '0' ELSE
      expandedKey_1(137);
  
  expandedKey_6(138) <= out0_112(138) WHEN out0_24 = '0' ELSE
      expandedKey_1(138);
  
  expandedKey_6(139) <= out0_112(139) WHEN out0_24 = '0' ELSE
      expandedKey_1(139);
  
  expandedKey_6(140) <= out0_112(140) WHEN out0_24 = '0' ELSE
      expandedKey_1(140);
  
  expandedKey_6(141) <= out0_112(141) WHEN out0_24 = '0' ELSE
      expandedKey_1(141);
  
  expandedKey_6(142) <= out0_112(142) WHEN out0_24 = '0' ELSE
      expandedKey_1(142);
  
  expandedKey_6(143) <= out0_112(143) WHEN out0_24 = '0' ELSE
      expandedKey_1(143);
  
  expandedKey_6(144) <= out0_112(144) WHEN out0_24 = '0' ELSE
      expandedKey_1(144);
  
  expandedKey_6(145) <= out0_112(145) WHEN out0_24 = '0' ELSE
      expandedKey_1(145);
  
  expandedKey_6(146) <= out0_112(146) WHEN out0_24 = '0' ELSE
      expandedKey_1(146);
  
  expandedKey_6(147) <= out0_112(147) WHEN out0_24 = '0' ELSE
      expandedKey_1(147);
  
  expandedKey_6(148) <= out0_112(148) WHEN out0_24 = '0' ELSE
      expandedKey_1(148);
  
  expandedKey_6(149) <= out0_112(149) WHEN out0_24 = '0' ELSE
      expandedKey_1(149);
  
  expandedKey_6(150) <= out0_112(150) WHEN out0_24 = '0' ELSE
      expandedKey_1(150);
  
  expandedKey_6(151) <= out0_112(151) WHEN out0_24 = '0' ELSE
      expandedKey_1(151);
  
  expandedKey_6(152) <= out0_112(152) WHEN out0_24 = '0' ELSE
      expandedKey_1(152);
  
  expandedKey_6(153) <= out0_112(153) WHEN out0_24 = '0' ELSE
      expandedKey_1(153);
  
  expandedKey_6(154) <= out0_112(154) WHEN out0_24 = '0' ELSE
      expandedKey_1(154);
  
  expandedKey_6(155) <= out0_112(155) WHEN out0_24 = '0' ELSE
      expandedKey_1(155);
  
  expandedKey_6(156) <= out0_112(156) WHEN out0_24 = '0' ELSE
      expandedKey_1(156);
  
  expandedKey_6(157) <= out0_112(157) WHEN out0_24 = '0' ELSE
      expandedKey_1(157);
  
  expandedKey_6(158) <= out0_112(158) WHEN out0_24 = '0' ELSE
      expandedKey_1(158);
  
  expandedKey_6(159) <= out0_112(159) WHEN out0_24 = '0' ELSE
      expandedKey_1(159);
  
  expandedKey_6(160) <= out0_112(160) WHEN out0_24 = '0' ELSE
      expandedKey_1(160);
  
  expandedKey_6(161) <= out0_112(161) WHEN out0_24 = '0' ELSE
      expandedKey_1(161);
  
  expandedKey_6(162) <= out0_112(162) WHEN out0_24 = '0' ELSE
      expandedKey_1(162);
  
  expandedKey_6(163) <= out0_112(163) WHEN out0_24 = '0' ELSE
      expandedKey_1(163);
  
  expandedKey_6(164) <= out0_112(164) WHEN out0_24 = '0' ELSE
      expandedKey_1(164);
  
  expandedKey_6(165) <= out0_112(165) WHEN out0_24 = '0' ELSE
      expandedKey_1(165);
  
  expandedKey_6(166) <= out0_112(166) WHEN out0_24 = '0' ELSE
      expandedKey_1(166);
  
  expandedKey_6(167) <= out0_112(167) WHEN out0_24 = '0' ELSE
      expandedKey_1(167);
  
  expandedKey_6(168) <= out0_112(168) WHEN out0_24 = '0' ELSE
      expandedKey_1(168);
  
  expandedKey_6(169) <= out0_112(169) WHEN out0_24 = '0' ELSE
      expandedKey_1(169);
  
  expandedKey_6(170) <= out0_112(170) WHEN out0_24 = '0' ELSE
      expandedKey_1(170);
  
  expandedKey_6(171) <= out0_112(171) WHEN out0_24 = '0' ELSE
      expandedKey_1(171);
  
  expandedKey_6(172) <= out0_112(172) WHEN out0_24 = '0' ELSE
      expandedKey_1(172);
  
  expandedKey_6(173) <= out0_112(173) WHEN out0_24 = '0' ELSE
      expandedKey_1(173);
  
  expandedKey_6(174) <= out0_112(174) WHEN out0_24 = '0' ELSE
      expandedKey_1(174);
  
  expandedKey_6(175) <= out0_112(175) WHEN out0_24 = '0' ELSE
      expandedKey_1(175);
  
  expandedKey_6(176) <= out0_112(176) WHEN out0_24 = '0' ELSE
      expandedKey_1(176);
  
  expandedKey_6(177) <= out0_112(177) WHEN out0_24 = '0' ELSE
      expandedKey_1(177);
  
  expandedKey_6(178) <= out0_112(178) WHEN out0_24 = '0' ELSE
      expandedKey_1(178);
  
  expandedKey_6(179) <= out0_112(179) WHEN out0_24 = '0' ELSE
      expandedKey_1(179);
  
  expandedKey_6(180) <= out0_112(180) WHEN out0_24 = '0' ELSE
      expandedKey_1(180);
  
  expandedKey_6(181) <= out0_112(181) WHEN out0_24 = '0' ELSE
      expandedKey_1(181);
  
  expandedKey_6(182) <= out0_112(182) WHEN out0_24 = '0' ELSE
      expandedKey_1(182);
  
  expandedKey_6(183) <= out0_112(183) WHEN out0_24 = '0' ELSE
      expandedKey_1(183);
  
  expandedKey_6(184) <= out0_112(184) WHEN out0_24 = '0' ELSE
      expandedKey_1(184);
  
  expandedKey_6(185) <= out0_112(185) WHEN out0_24 = '0' ELSE
      expandedKey_1(185);
  
  expandedKey_6(186) <= out0_112(186) WHEN out0_24 = '0' ELSE
      expandedKey_1(186);
  
  expandedKey_6(187) <= out0_112(187) WHEN out0_24 = '0' ELSE
      expandedKey_1(187);
  
  expandedKey_6(188) <= out0_112(188) WHEN out0_24 = '0' ELSE
      expandedKey_1(188);
  
  expandedKey_6(189) <= out0_112(189) WHEN out0_24 = '0' ELSE
      expandedKey_1(189);
  
  expandedKey_6(190) <= out0_112(190) WHEN out0_24 = '0' ELSE
      expandedKey_1(190);
  
  expandedKey_6(191) <= out0_112(191) WHEN out0_24 = '0' ELSE
      expandedKey_1(191);
  
  expandedKey_6(192) <= out0_112(192) WHEN out0_24 = '0' ELSE
      expandedKey_1(192);
  
  expandedKey_6(193) <= out0_112(193) WHEN out0_24 = '0' ELSE
      expandedKey_1(193);
  
  expandedKey_6(194) <= out0_112(194) WHEN out0_24 = '0' ELSE
      expandedKey_1(194);
  
  expandedKey_6(195) <= out0_112(195) WHEN out0_24 = '0' ELSE
      expandedKey_1(195);
  
  expandedKey_6(196) <= out0_112(196) WHEN out0_24 = '0' ELSE
      expandedKey_1(196);
  
  expandedKey_6(197) <= out0_112(197) WHEN out0_24 = '0' ELSE
      expandedKey_1(197);
  
  expandedKey_6(198) <= out0_112(198) WHEN out0_24 = '0' ELSE
      expandedKey_1(198);
  
  expandedKey_6(199) <= out0_112(199) WHEN out0_24 = '0' ELSE
      expandedKey_1(199);
  
  expandedKey_6(200) <= out0_112(200) WHEN out0_24 = '0' ELSE
      expandedKey_1(200);
  
  expandedKey_6(201) <= out0_112(201) WHEN out0_24 = '0' ELSE
      expandedKey_1(201);
  
  expandedKey_6(202) <= out0_112(202) WHEN out0_24 = '0' ELSE
      expandedKey_1(202);
  
  expandedKey_6(203) <= out0_112(203) WHEN out0_24 = '0' ELSE
      expandedKey_1(203);
  
  expandedKey_6(204) <= out0_112(204) WHEN out0_24 = '0' ELSE
      expandedKey_1(204);
  
  expandedKey_6(205) <= out0_112(205) WHEN out0_24 = '0' ELSE
      expandedKey_1(205);
  
  expandedKey_6(206) <= out0_112(206) WHEN out0_24 = '0' ELSE
      expandedKey_1(206);
  
  expandedKey_6(207) <= out0_112(207) WHEN out0_24 = '0' ELSE
      expandedKey_1(207);
  
  expandedKey_6(208) <= out0_112(208) WHEN out0_24 = '0' ELSE
      expandedKey_1(208);
  
  expandedKey_6(209) <= out0_112(209) WHEN out0_24 = '0' ELSE
      expandedKey_1(209);
  
  expandedKey_6(210) <= out0_112(210) WHEN out0_24 = '0' ELSE
      expandedKey_1(210);
  
  expandedKey_6(211) <= out0_112(211) WHEN out0_24 = '0' ELSE
      expandedKey_1(211);
  
  expandedKey_6(212) <= out0_112(212) WHEN out0_24 = '0' ELSE
      expandedKey_1(212);
  
  expandedKey_6(213) <= out0_112(213) WHEN out0_24 = '0' ELSE
      expandedKey_1(213);
  
  expandedKey_6(214) <= out0_112(214) WHEN out0_24 = '0' ELSE
      expandedKey_1(214);
  
  expandedKey_6(215) <= out0_112(215) WHEN out0_24 = '0' ELSE
      expandedKey_1(215);
  
  expandedKey_6(216) <= out0_112(216) WHEN out0_24 = '0' ELSE
      expandedKey_1(216);
  
  expandedKey_6(217) <= out0_112(217) WHEN out0_24 = '0' ELSE
      expandedKey_1(217);
  
  expandedKey_6(218) <= out0_112(218) WHEN out0_24 = '0' ELSE
      expandedKey_1(218);
  
  expandedKey_6(219) <= out0_112(219) WHEN out0_24 = '0' ELSE
      expandedKey_1(219);
  
  expandedKey_6(220) <= out0_112(220) WHEN out0_24 = '0' ELSE
      expandedKey_1(220);
  
  expandedKey_6(221) <= out0_112(221) WHEN out0_24 = '0' ELSE
      expandedKey_1(221);
  
  expandedKey_6(222) <= out0_112(222) WHEN out0_24 = '0' ELSE
      expandedKey_1(222);
  
  expandedKey_6(223) <= out0_112(223) WHEN out0_24 = '0' ELSE
      expandedKey_1(223);
  
  expandedKey_6(224) <= out0_112(224) WHEN out0_24 = '0' ELSE
      expandedKey_1(224);
  
  expandedKey_6(225) <= out0_112(225) WHEN out0_24 = '0' ELSE
      expandedKey_1(225);
  
  expandedKey_6(226) <= out0_112(226) WHEN out0_24 = '0' ELSE
      expandedKey_1(226);
  
  expandedKey_6(227) <= out0_112(227) WHEN out0_24 = '0' ELSE
      expandedKey_1(227);
  
  expandedKey_6(228) <= out0_112(228) WHEN out0_24 = '0' ELSE
      expandedKey_1(228);
  
  expandedKey_6(229) <= out0_112(229) WHEN out0_24 = '0' ELSE
      expandedKey_1(229);
  
  expandedKey_6(230) <= out0_112(230) WHEN out0_24 = '0' ELSE
      expandedKey_1(230);
  
  expandedKey_6(231) <= out0_112(231) WHEN out0_24 = '0' ELSE
      expandedKey_1(231);
  
  expandedKey_6(232) <= out0_112(232) WHEN out0_24 = '0' ELSE
      expandedKey_1(232);
  
  expandedKey_6(233) <= out0_112(233) WHEN out0_24 = '0' ELSE
      expandedKey_1(233);
  
  expandedKey_6(234) <= out0_112(234) WHEN out0_24 = '0' ELSE
      expandedKey_1(234);
  
  expandedKey_6(235) <= out0_112(235) WHEN out0_24 = '0' ELSE
      expandedKey_1(235);
  
  expandedKey_6(236) <= out0_112(236) WHEN out0_24 = '0' ELSE
      expandedKey_1(236);
  
  expandedKey_6(237) <= out0_112(237) WHEN out0_24 = '0' ELSE
      expandedKey_1(237);
  
  expandedKey_6(238) <= out0_112(238) WHEN out0_24 = '0' ELSE
      expandedKey_1(238);
  
  expandedKey_6(239) <= out0_112(239) WHEN out0_24 = '0' ELSE
      expandedKey_1(239);

  intdelay5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        expandedKey(0) <= to_unsigned(16#00#, 8);
        expandedKey(1) <= to_unsigned(16#00#, 8);
        expandedKey(2) <= to_unsigned(16#00#, 8);
        expandedKey(3) <= to_unsigned(16#00#, 8);
        expandedKey(4) <= to_unsigned(16#00#, 8);
        expandedKey(5) <= to_unsigned(16#00#, 8);
        expandedKey(6) <= to_unsigned(16#00#, 8);
        expandedKey(7) <= to_unsigned(16#00#, 8);
        expandedKey(8) <= to_unsigned(16#00#, 8);
        expandedKey(9) <= to_unsigned(16#00#, 8);
        expandedKey(10) <= to_unsigned(16#00#, 8);
        expandedKey(11) <= to_unsigned(16#00#, 8);
        expandedKey(12) <= to_unsigned(16#00#, 8);
        expandedKey(13) <= to_unsigned(16#00#, 8);
        expandedKey(14) <= to_unsigned(16#00#, 8);
        expandedKey(15) <= to_unsigned(16#00#, 8);
        expandedKey(16) <= to_unsigned(16#00#, 8);
        expandedKey(17) <= to_unsigned(16#00#, 8);
        expandedKey(18) <= to_unsigned(16#00#, 8);
        expandedKey(19) <= to_unsigned(16#00#, 8);
        expandedKey(20) <= to_unsigned(16#00#, 8);
        expandedKey(21) <= to_unsigned(16#00#, 8);
        expandedKey(22) <= to_unsigned(16#00#, 8);
        expandedKey(23) <= to_unsigned(16#00#, 8);
        expandedKey(24) <= to_unsigned(16#00#, 8);
        expandedKey(25) <= to_unsigned(16#00#, 8);
        expandedKey(26) <= to_unsigned(16#00#, 8);
        expandedKey(27) <= to_unsigned(16#00#, 8);
        expandedKey(28) <= to_unsigned(16#00#, 8);
        expandedKey(29) <= to_unsigned(16#00#, 8);
        expandedKey(30) <= to_unsigned(16#00#, 8);
        expandedKey(31) <= to_unsigned(16#00#, 8);
        expandedKey(32) <= to_unsigned(16#00#, 8);
        expandedKey(33) <= to_unsigned(16#00#, 8);
        expandedKey(34) <= to_unsigned(16#00#, 8);
        expandedKey(35) <= to_unsigned(16#00#, 8);
        expandedKey(36) <= to_unsigned(16#00#, 8);
        expandedKey(37) <= to_unsigned(16#00#, 8);
        expandedKey(38) <= to_unsigned(16#00#, 8);
        expandedKey(39) <= to_unsigned(16#00#, 8);
        expandedKey(40) <= to_unsigned(16#00#, 8);
        expandedKey(41) <= to_unsigned(16#00#, 8);
        expandedKey(42) <= to_unsigned(16#00#, 8);
        expandedKey(43) <= to_unsigned(16#00#, 8);
        expandedKey(44) <= to_unsigned(16#00#, 8);
        expandedKey(45) <= to_unsigned(16#00#, 8);
        expandedKey(46) <= to_unsigned(16#00#, 8);
        expandedKey(47) <= to_unsigned(16#00#, 8);
        expandedKey(48) <= to_unsigned(16#00#, 8);
        expandedKey(49) <= to_unsigned(16#00#, 8);
        expandedKey(50) <= to_unsigned(16#00#, 8);
        expandedKey(51) <= to_unsigned(16#00#, 8);
        expandedKey(52) <= to_unsigned(16#00#, 8);
        expandedKey(53) <= to_unsigned(16#00#, 8);
        expandedKey(54) <= to_unsigned(16#00#, 8);
        expandedKey(55) <= to_unsigned(16#00#, 8);
        expandedKey(56) <= to_unsigned(16#00#, 8);
        expandedKey(57) <= to_unsigned(16#00#, 8);
        expandedKey(58) <= to_unsigned(16#00#, 8);
        expandedKey(59) <= to_unsigned(16#00#, 8);
        expandedKey(60) <= to_unsigned(16#00#, 8);
        expandedKey(61) <= to_unsigned(16#00#, 8);
        expandedKey(62) <= to_unsigned(16#00#, 8);
        expandedKey(63) <= to_unsigned(16#00#, 8);
        expandedKey(64) <= to_unsigned(16#00#, 8);
        expandedKey(65) <= to_unsigned(16#00#, 8);
        expandedKey(66) <= to_unsigned(16#00#, 8);
        expandedKey(67) <= to_unsigned(16#00#, 8);
        expandedKey(68) <= to_unsigned(16#00#, 8);
        expandedKey(69) <= to_unsigned(16#00#, 8);
        expandedKey(70) <= to_unsigned(16#00#, 8);
        expandedKey(71) <= to_unsigned(16#00#, 8);
        expandedKey(72) <= to_unsigned(16#00#, 8);
        expandedKey(73) <= to_unsigned(16#00#, 8);
        expandedKey(74) <= to_unsigned(16#00#, 8);
        expandedKey(75) <= to_unsigned(16#00#, 8);
        expandedKey(76) <= to_unsigned(16#00#, 8);
        expandedKey(77) <= to_unsigned(16#00#, 8);
        expandedKey(78) <= to_unsigned(16#00#, 8);
        expandedKey(79) <= to_unsigned(16#00#, 8);
        expandedKey(80) <= to_unsigned(16#00#, 8);
        expandedKey(81) <= to_unsigned(16#00#, 8);
        expandedKey(82) <= to_unsigned(16#00#, 8);
        expandedKey(83) <= to_unsigned(16#00#, 8);
        expandedKey(84) <= to_unsigned(16#00#, 8);
        expandedKey(85) <= to_unsigned(16#00#, 8);
        expandedKey(86) <= to_unsigned(16#00#, 8);
        expandedKey(87) <= to_unsigned(16#00#, 8);
        expandedKey(88) <= to_unsigned(16#00#, 8);
        expandedKey(89) <= to_unsigned(16#00#, 8);
        expandedKey(90) <= to_unsigned(16#00#, 8);
        expandedKey(91) <= to_unsigned(16#00#, 8);
        expandedKey(92) <= to_unsigned(16#00#, 8);
        expandedKey(93) <= to_unsigned(16#00#, 8);
        expandedKey(94) <= to_unsigned(16#00#, 8);
        expandedKey(95) <= to_unsigned(16#00#, 8);
        expandedKey(96) <= to_unsigned(16#00#, 8);
        expandedKey(97) <= to_unsigned(16#00#, 8);
        expandedKey(98) <= to_unsigned(16#00#, 8);
        expandedKey(99) <= to_unsigned(16#00#, 8);
        expandedKey(100) <= to_unsigned(16#00#, 8);
        expandedKey(101) <= to_unsigned(16#00#, 8);
        expandedKey(102) <= to_unsigned(16#00#, 8);
        expandedKey(103) <= to_unsigned(16#00#, 8);
        expandedKey(104) <= to_unsigned(16#00#, 8);
        expandedKey(105) <= to_unsigned(16#00#, 8);
        expandedKey(106) <= to_unsigned(16#00#, 8);
        expandedKey(107) <= to_unsigned(16#00#, 8);
        expandedKey(108) <= to_unsigned(16#00#, 8);
        expandedKey(109) <= to_unsigned(16#00#, 8);
        expandedKey(110) <= to_unsigned(16#00#, 8);
        expandedKey(111) <= to_unsigned(16#00#, 8);
        expandedKey(112) <= to_unsigned(16#00#, 8);
        expandedKey(113) <= to_unsigned(16#00#, 8);
        expandedKey(114) <= to_unsigned(16#00#, 8);
        expandedKey(115) <= to_unsigned(16#00#, 8);
        expandedKey(116) <= to_unsigned(16#00#, 8);
        expandedKey(117) <= to_unsigned(16#00#, 8);
        expandedKey(118) <= to_unsigned(16#00#, 8);
        expandedKey(119) <= to_unsigned(16#00#, 8);
        expandedKey(120) <= to_unsigned(16#00#, 8);
        expandedKey(121) <= to_unsigned(16#00#, 8);
        expandedKey(122) <= to_unsigned(16#00#, 8);
        expandedKey(123) <= to_unsigned(16#00#, 8);
        expandedKey(124) <= to_unsigned(16#00#, 8);
        expandedKey(125) <= to_unsigned(16#00#, 8);
        expandedKey(126) <= to_unsigned(16#00#, 8);
        expandedKey(127) <= to_unsigned(16#00#, 8);
        expandedKey(128) <= to_unsigned(16#00#, 8);
        expandedKey(129) <= to_unsigned(16#00#, 8);
        expandedKey(130) <= to_unsigned(16#00#, 8);
        expandedKey(131) <= to_unsigned(16#00#, 8);
        expandedKey(132) <= to_unsigned(16#00#, 8);
        expandedKey(133) <= to_unsigned(16#00#, 8);
        expandedKey(134) <= to_unsigned(16#00#, 8);
        expandedKey(135) <= to_unsigned(16#00#, 8);
        expandedKey(136) <= to_unsigned(16#00#, 8);
        expandedKey(137) <= to_unsigned(16#00#, 8);
        expandedKey(138) <= to_unsigned(16#00#, 8);
        expandedKey(139) <= to_unsigned(16#00#, 8);
        expandedKey(140) <= to_unsigned(16#00#, 8);
        expandedKey(141) <= to_unsigned(16#00#, 8);
        expandedKey(142) <= to_unsigned(16#00#, 8);
        expandedKey(143) <= to_unsigned(16#00#, 8);
        expandedKey(144) <= to_unsigned(16#00#, 8);
        expandedKey(145) <= to_unsigned(16#00#, 8);
        expandedKey(146) <= to_unsigned(16#00#, 8);
        expandedKey(147) <= to_unsigned(16#00#, 8);
        expandedKey(148) <= to_unsigned(16#00#, 8);
        expandedKey(149) <= to_unsigned(16#00#, 8);
        expandedKey(150) <= to_unsigned(16#00#, 8);
        expandedKey(151) <= to_unsigned(16#00#, 8);
        expandedKey(152) <= to_unsigned(16#00#, 8);
        expandedKey(153) <= to_unsigned(16#00#, 8);
        expandedKey(154) <= to_unsigned(16#00#, 8);
        expandedKey(155) <= to_unsigned(16#00#, 8);
        expandedKey(156) <= to_unsigned(16#00#, 8);
        expandedKey(157) <= to_unsigned(16#00#, 8);
        expandedKey(158) <= to_unsigned(16#00#, 8);
        expandedKey(159) <= to_unsigned(16#00#, 8);
        expandedKey(160) <= to_unsigned(16#00#, 8);
        expandedKey(161) <= to_unsigned(16#00#, 8);
        expandedKey(162) <= to_unsigned(16#00#, 8);
        expandedKey(163) <= to_unsigned(16#00#, 8);
        expandedKey(164) <= to_unsigned(16#00#, 8);
        expandedKey(165) <= to_unsigned(16#00#, 8);
        expandedKey(166) <= to_unsigned(16#00#, 8);
        expandedKey(167) <= to_unsigned(16#00#, 8);
        expandedKey(168) <= to_unsigned(16#00#, 8);
        expandedKey(169) <= to_unsigned(16#00#, 8);
        expandedKey(170) <= to_unsigned(16#00#, 8);
        expandedKey(171) <= to_unsigned(16#00#, 8);
        expandedKey(172) <= to_unsigned(16#00#, 8);
        expandedKey(173) <= to_unsigned(16#00#, 8);
        expandedKey(174) <= to_unsigned(16#00#, 8);
        expandedKey(175) <= to_unsigned(16#00#, 8);
        expandedKey(176) <= to_unsigned(16#00#, 8);
        expandedKey(177) <= to_unsigned(16#00#, 8);
        expandedKey(178) <= to_unsigned(16#00#, 8);
        expandedKey(179) <= to_unsigned(16#00#, 8);
        expandedKey(180) <= to_unsigned(16#00#, 8);
        expandedKey(181) <= to_unsigned(16#00#, 8);
        expandedKey(182) <= to_unsigned(16#00#, 8);
        expandedKey(183) <= to_unsigned(16#00#, 8);
        expandedKey(184) <= to_unsigned(16#00#, 8);
        expandedKey(185) <= to_unsigned(16#00#, 8);
        expandedKey(186) <= to_unsigned(16#00#, 8);
        expandedKey(187) <= to_unsigned(16#00#, 8);
        expandedKey(188) <= to_unsigned(16#00#, 8);
        expandedKey(189) <= to_unsigned(16#00#, 8);
        expandedKey(190) <= to_unsigned(16#00#, 8);
        expandedKey(191) <= to_unsigned(16#00#, 8);
        expandedKey(192) <= to_unsigned(16#00#, 8);
        expandedKey(193) <= to_unsigned(16#00#, 8);
        expandedKey(194) <= to_unsigned(16#00#, 8);
        expandedKey(195) <= to_unsigned(16#00#, 8);
        expandedKey(196) <= to_unsigned(16#00#, 8);
        expandedKey(197) <= to_unsigned(16#00#, 8);
        expandedKey(198) <= to_unsigned(16#00#, 8);
        expandedKey(199) <= to_unsigned(16#00#, 8);
        expandedKey(200) <= to_unsigned(16#00#, 8);
        expandedKey(201) <= to_unsigned(16#00#, 8);
        expandedKey(202) <= to_unsigned(16#00#, 8);
        expandedKey(203) <= to_unsigned(16#00#, 8);
        expandedKey(204) <= to_unsigned(16#00#, 8);
        expandedKey(205) <= to_unsigned(16#00#, 8);
        expandedKey(206) <= to_unsigned(16#00#, 8);
        expandedKey(207) <= to_unsigned(16#00#, 8);
        expandedKey(208) <= to_unsigned(16#00#, 8);
        expandedKey(209) <= to_unsigned(16#00#, 8);
        expandedKey(210) <= to_unsigned(16#00#, 8);
        expandedKey(211) <= to_unsigned(16#00#, 8);
        expandedKey(212) <= to_unsigned(16#00#, 8);
        expandedKey(213) <= to_unsigned(16#00#, 8);
        expandedKey(214) <= to_unsigned(16#00#, 8);
        expandedKey(215) <= to_unsigned(16#00#, 8);
        expandedKey(216) <= to_unsigned(16#00#, 8);
        expandedKey(217) <= to_unsigned(16#00#, 8);
        expandedKey(218) <= to_unsigned(16#00#, 8);
        expandedKey(219) <= to_unsigned(16#00#, 8);
        expandedKey(220) <= to_unsigned(16#00#, 8);
        expandedKey(221) <= to_unsigned(16#00#, 8);
        expandedKey(222) <= to_unsigned(16#00#, 8);
        expandedKey(223) <= to_unsigned(16#00#, 8);
        expandedKey(224) <= to_unsigned(16#00#, 8);
        expandedKey(225) <= to_unsigned(16#00#, 8);
        expandedKey(226) <= to_unsigned(16#00#, 8);
        expandedKey(227) <= to_unsigned(16#00#, 8);
        expandedKey(228) <= to_unsigned(16#00#, 8);
        expandedKey(229) <= to_unsigned(16#00#, 8);
        expandedKey(230) <= to_unsigned(16#00#, 8);
        expandedKey(231) <= to_unsigned(16#00#, 8);
        expandedKey(232) <= to_unsigned(16#00#, 8);
        expandedKey(233) <= to_unsigned(16#00#, 8);
        expandedKey(234) <= to_unsigned(16#00#, 8);
        expandedKey(235) <= to_unsigned(16#00#, 8);
        expandedKey(236) <= to_unsigned(16#00#, 8);
        expandedKey(237) <= to_unsigned(16#00#, 8);
        expandedKey(238) <= to_unsigned(16#00#, 8);
        expandedKey(239) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        expandedKey(0) <= expandedKey_6(0);
        expandedKey(1) <= expandedKey_6(1);
        expandedKey(2) <= expandedKey_6(2);
        expandedKey(3) <= expandedKey_6(3);
        expandedKey(4) <= expandedKey_6(4);
        expandedKey(5) <= expandedKey_6(5);
        expandedKey(6) <= expandedKey_6(6);
        expandedKey(7) <= expandedKey_6(7);
        expandedKey(8) <= expandedKey_6(8);
        expandedKey(9) <= expandedKey_6(9);
        expandedKey(10) <= expandedKey_6(10);
        expandedKey(11) <= expandedKey_6(11);
        expandedKey(12) <= expandedKey_6(12);
        expandedKey(13) <= expandedKey_6(13);
        expandedKey(14) <= expandedKey_6(14);
        expandedKey(15) <= expandedKey_6(15);
        expandedKey(16) <= expandedKey_6(16);
        expandedKey(17) <= expandedKey_6(17);
        expandedKey(18) <= expandedKey_6(18);
        expandedKey(19) <= expandedKey_6(19);
        expandedKey(20) <= expandedKey_6(20);
        expandedKey(21) <= expandedKey_6(21);
        expandedKey(22) <= expandedKey_6(22);
        expandedKey(23) <= expandedKey_6(23);
        expandedKey(24) <= expandedKey_6(24);
        expandedKey(25) <= expandedKey_6(25);
        expandedKey(26) <= expandedKey_6(26);
        expandedKey(27) <= expandedKey_6(27);
        expandedKey(28) <= expandedKey_6(28);
        expandedKey(29) <= expandedKey_6(29);
        expandedKey(30) <= expandedKey_6(30);
        expandedKey(31) <= expandedKey_6(31);
        expandedKey(32) <= expandedKey_6(32);
        expandedKey(33) <= expandedKey_6(33);
        expandedKey(34) <= expandedKey_6(34);
        expandedKey(35) <= expandedKey_6(35);
        expandedKey(36) <= expandedKey_6(36);
        expandedKey(37) <= expandedKey_6(37);
        expandedKey(38) <= expandedKey_6(38);
        expandedKey(39) <= expandedKey_6(39);
        expandedKey(40) <= expandedKey_6(40);
        expandedKey(41) <= expandedKey_6(41);
        expandedKey(42) <= expandedKey_6(42);
        expandedKey(43) <= expandedKey_6(43);
        expandedKey(44) <= expandedKey_6(44);
        expandedKey(45) <= expandedKey_6(45);
        expandedKey(46) <= expandedKey_6(46);
        expandedKey(47) <= expandedKey_6(47);
        expandedKey(48) <= expandedKey_6(48);
        expandedKey(49) <= expandedKey_6(49);
        expandedKey(50) <= expandedKey_6(50);
        expandedKey(51) <= expandedKey_6(51);
        expandedKey(52) <= expandedKey_6(52);
        expandedKey(53) <= expandedKey_6(53);
        expandedKey(54) <= expandedKey_6(54);
        expandedKey(55) <= expandedKey_6(55);
        expandedKey(56) <= expandedKey_6(56);
        expandedKey(57) <= expandedKey_6(57);
        expandedKey(58) <= expandedKey_6(58);
        expandedKey(59) <= expandedKey_6(59);
        expandedKey(60) <= expandedKey_6(60);
        expandedKey(61) <= expandedKey_6(61);
        expandedKey(62) <= expandedKey_6(62);
        expandedKey(63) <= expandedKey_6(63);
        expandedKey(64) <= expandedKey_6(64);
        expandedKey(65) <= expandedKey_6(65);
        expandedKey(66) <= expandedKey_6(66);
        expandedKey(67) <= expandedKey_6(67);
        expandedKey(68) <= expandedKey_6(68);
        expandedKey(69) <= expandedKey_6(69);
        expandedKey(70) <= expandedKey_6(70);
        expandedKey(71) <= expandedKey_6(71);
        expandedKey(72) <= expandedKey_6(72);
        expandedKey(73) <= expandedKey_6(73);
        expandedKey(74) <= expandedKey_6(74);
        expandedKey(75) <= expandedKey_6(75);
        expandedKey(76) <= expandedKey_6(76);
        expandedKey(77) <= expandedKey_6(77);
        expandedKey(78) <= expandedKey_6(78);
        expandedKey(79) <= expandedKey_6(79);
        expandedKey(80) <= expandedKey_6(80);
        expandedKey(81) <= expandedKey_6(81);
        expandedKey(82) <= expandedKey_6(82);
        expandedKey(83) <= expandedKey_6(83);
        expandedKey(84) <= expandedKey_6(84);
        expandedKey(85) <= expandedKey_6(85);
        expandedKey(86) <= expandedKey_6(86);
        expandedKey(87) <= expandedKey_6(87);
        expandedKey(88) <= expandedKey_6(88);
        expandedKey(89) <= expandedKey_6(89);
        expandedKey(90) <= expandedKey_6(90);
        expandedKey(91) <= expandedKey_6(91);
        expandedKey(92) <= expandedKey_6(92);
        expandedKey(93) <= expandedKey_6(93);
        expandedKey(94) <= expandedKey_6(94);
        expandedKey(95) <= expandedKey_6(95);
        expandedKey(96) <= expandedKey_6(96);
        expandedKey(97) <= expandedKey_6(97);
        expandedKey(98) <= expandedKey_6(98);
        expandedKey(99) <= expandedKey_6(99);
        expandedKey(100) <= expandedKey_6(100);
        expandedKey(101) <= expandedKey_6(101);
        expandedKey(102) <= expandedKey_6(102);
        expandedKey(103) <= expandedKey_6(103);
        expandedKey(104) <= expandedKey_6(104);
        expandedKey(105) <= expandedKey_6(105);
        expandedKey(106) <= expandedKey_6(106);
        expandedKey(107) <= expandedKey_6(107);
        expandedKey(108) <= expandedKey_6(108);
        expandedKey(109) <= expandedKey_6(109);
        expandedKey(110) <= expandedKey_6(110);
        expandedKey(111) <= expandedKey_6(111);
        expandedKey(112) <= expandedKey_6(112);
        expandedKey(113) <= expandedKey_6(113);
        expandedKey(114) <= expandedKey_6(114);
        expandedKey(115) <= expandedKey_6(115);
        expandedKey(116) <= expandedKey_6(116);
        expandedKey(117) <= expandedKey_6(117);
        expandedKey(118) <= expandedKey_6(118);
        expandedKey(119) <= expandedKey_6(119);
        expandedKey(120) <= expandedKey_6(120);
        expandedKey(121) <= expandedKey_6(121);
        expandedKey(122) <= expandedKey_6(122);
        expandedKey(123) <= expandedKey_6(123);
        expandedKey(124) <= expandedKey_6(124);
        expandedKey(125) <= expandedKey_6(125);
        expandedKey(126) <= expandedKey_6(126);
        expandedKey(127) <= expandedKey_6(127);
        expandedKey(128) <= expandedKey_6(128);
        expandedKey(129) <= expandedKey_6(129);
        expandedKey(130) <= expandedKey_6(130);
        expandedKey(131) <= expandedKey_6(131);
        expandedKey(132) <= expandedKey_6(132);
        expandedKey(133) <= expandedKey_6(133);
        expandedKey(134) <= expandedKey_6(134);
        expandedKey(135) <= expandedKey_6(135);
        expandedKey(136) <= expandedKey_6(136);
        expandedKey(137) <= expandedKey_6(137);
        expandedKey(138) <= expandedKey_6(138);
        expandedKey(139) <= expandedKey_6(139);
        expandedKey(140) <= expandedKey_6(140);
        expandedKey(141) <= expandedKey_6(141);
        expandedKey(142) <= expandedKey_6(142);
        expandedKey(143) <= expandedKey_6(143);
        expandedKey(144) <= expandedKey_6(144);
        expandedKey(145) <= expandedKey_6(145);
        expandedKey(146) <= expandedKey_6(146);
        expandedKey(147) <= expandedKey_6(147);
        expandedKey(148) <= expandedKey_6(148);
        expandedKey(149) <= expandedKey_6(149);
        expandedKey(150) <= expandedKey_6(150);
        expandedKey(151) <= expandedKey_6(151);
        expandedKey(152) <= expandedKey_6(152);
        expandedKey(153) <= expandedKey_6(153);
        expandedKey(154) <= expandedKey_6(154);
        expandedKey(155) <= expandedKey_6(155);
        expandedKey(156) <= expandedKey_6(156);
        expandedKey(157) <= expandedKey_6(157);
        expandedKey(158) <= expandedKey_6(158);
        expandedKey(159) <= expandedKey_6(159);
        expandedKey(160) <= expandedKey_6(160);
        expandedKey(161) <= expandedKey_6(161);
        expandedKey(162) <= expandedKey_6(162);
        expandedKey(163) <= expandedKey_6(163);
        expandedKey(164) <= expandedKey_6(164);
        expandedKey(165) <= expandedKey_6(165);
        expandedKey(166) <= expandedKey_6(166);
        expandedKey(167) <= expandedKey_6(167);
        expandedKey(168) <= expandedKey_6(168);
        expandedKey(169) <= expandedKey_6(169);
        expandedKey(170) <= expandedKey_6(170);
        expandedKey(171) <= expandedKey_6(171);
        expandedKey(172) <= expandedKey_6(172);
        expandedKey(173) <= expandedKey_6(173);
        expandedKey(174) <= expandedKey_6(174);
        expandedKey(175) <= expandedKey_6(175);
        expandedKey(176) <= expandedKey_6(176);
        expandedKey(177) <= expandedKey_6(177);
        expandedKey(178) <= expandedKey_6(178);
        expandedKey(179) <= expandedKey_6(179);
        expandedKey(180) <= expandedKey_6(180);
        expandedKey(181) <= expandedKey_6(181);
        expandedKey(182) <= expandedKey_6(182);
        expandedKey(183) <= expandedKey_6(183);
        expandedKey(184) <= expandedKey_6(184);
        expandedKey(185) <= expandedKey_6(185);
        expandedKey(186) <= expandedKey_6(186);
        expandedKey(187) <= expandedKey_6(187);
        expandedKey(188) <= expandedKey_6(188);
        expandedKey(189) <= expandedKey_6(189);
        expandedKey(190) <= expandedKey_6(190);
        expandedKey(191) <= expandedKey_6(191);
        expandedKey(192) <= expandedKey_6(192);
        expandedKey(193) <= expandedKey_6(193);
        expandedKey(194) <= expandedKey_6(194);
        expandedKey(195) <= expandedKey_6(195);
        expandedKey(196) <= expandedKey_6(196);
        expandedKey(197) <= expandedKey_6(197);
        expandedKey(198) <= expandedKey_6(198);
        expandedKey(199) <= expandedKey_6(199);
        expandedKey(200) <= expandedKey_6(200);
        expandedKey(201) <= expandedKey_6(201);
        expandedKey(202) <= expandedKey_6(202);
        expandedKey(203) <= expandedKey_6(203);
        expandedKey(204) <= expandedKey_6(204);
        expandedKey(205) <= expandedKey_6(205);
        expandedKey(206) <= expandedKey_6(206);
        expandedKey(207) <= expandedKey_6(207);
        expandedKey(208) <= expandedKey_6(208);
        expandedKey(209) <= expandedKey_6(209);
        expandedKey(210) <= expandedKey_6(210);
        expandedKey(211) <= expandedKey_6(211);
        expandedKey(212) <= expandedKey_6(212);
        expandedKey(213) <= expandedKey_6(213);
        expandedKey(214) <= expandedKey_6(214);
        expandedKey(215) <= expandedKey_6(215);
        expandedKey(216) <= expandedKey_6(216);
        expandedKey(217) <= expandedKey_6(217);
        expandedKey(218) <= expandedKey_6(218);
        expandedKey(219) <= expandedKey_6(219);
        expandedKey(220) <= expandedKey_6(220);
        expandedKey(221) <= expandedKey_6(221);
        expandedKey(222) <= expandedKey_6(222);
        expandedKey(223) <= expandedKey_6(223);
        expandedKey(224) <= expandedKey_6(224);
        expandedKey(225) <= expandedKey_6(225);
        expandedKey(226) <= expandedKey_6(226);
        expandedKey(227) <= expandedKey_6(227);
        expandedKey(228) <= expandedKey_6(228);
        expandedKey(229) <= expandedKey_6(229);
        expandedKey(230) <= expandedKey_6(230);
        expandedKey(231) <= expandedKey_6(231);
        expandedKey(232) <= expandedKey_6(232);
        expandedKey(233) <= expandedKey_6(233);
        expandedKey(234) <= expandedKey_6(234);
        expandedKey(235) <= expandedKey_6(235);
        expandedKey(236) <= expandedKey_6(236);
        expandedKey(237) <= expandedKey_6(237);
        expandedKey(238) <= expandedKey_6(238);
        expandedKey(239) <= expandedKey_6(239);
      END IF;
    END IF;
  END PROCESS intdelay5_process;


  
  out0_113 <= expandedKey(0) WHEN out0_49 = to_unsigned(16#01#, 8) ELSE
      expandedKey(1) WHEN out0_49 = to_unsigned(16#02#, 8) ELSE
      expandedKey(2) WHEN out0_49 = to_unsigned(16#03#, 8) ELSE
      expandedKey(3) WHEN out0_49 = to_unsigned(16#04#, 8) ELSE
      expandedKey(4) WHEN out0_49 = to_unsigned(16#05#, 8) ELSE
      expandedKey(5) WHEN out0_49 = to_unsigned(16#06#, 8) ELSE
      expandedKey(6) WHEN out0_49 = to_unsigned(16#07#, 8) ELSE
      expandedKey(7) WHEN out0_49 = to_unsigned(16#08#, 8) ELSE
      expandedKey(8) WHEN out0_49 = to_unsigned(16#09#, 8) ELSE
      expandedKey(9) WHEN out0_49 = to_unsigned(16#0A#, 8) ELSE
      expandedKey(10) WHEN out0_49 = to_unsigned(16#0B#, 8) ELSE
      expandedKey(11) WHEN out0_49 = to_unsigned(16#0C#, 8) ELSE
      expandedKey(12) WHEN out0_49 = to_unsigned(16#0D#, 8) ELSE
      expandedKey(13) WHEN out0_49 = to_unsigned(16#0E#, 8) ELSE
      expandedKey(14) WHEN out0_49 = to_unsigned(16#0F#, 8) ELSE
      expandedKey(15) WHEN out0_49 = to_unsigned(16#10#, 8) ELSE
      expandedKey(16) WHEN out0_49 = to_unsigned(16#11#, 8) ELSE
      expandedKey(17) WHEN out0_49 = to_unsigned(16#12#, 8) ELSE
      expandedKey(18) WHEN out0_49 = to_unsigned(16#13#, 8) ELSE
      expandedKey(19) WHEN out0_49 = to_unsigned(16#14#, 8) ELSE
      expandedKey(20) WHEN out0_49 = to_unsigned(16#15#, 8) ELSE
      expandedKey(21) WHEN out0_49 = to_unsigned(16#16#, 8) ELSE
      expandedKey(22) WHEN out0_49 = to_unsigned(16#17#, 8) ELSE
      expandedKey(23) WHEN out0_49 = to_unsigned(16#18#, 8) ELSE
      expandedKey(24) WHEN out0_49 = to_unsigned(16#19#, 8) ELSE
      expandedKey(25) WHEN out0_49 = to_unsigned(16#1A#, 8) ELSE
      expandedKey(26) WHEN out0_49 = to_unsigned(16#1B#, 8) ELSE
      expandedKey(27) WHEN out0_49 = to_unsigned(16#1C#, 8) ELSE
      expandedKey(28) WHEN out0_49 = to_unsigned(16#1D#, 8) ELSE
      expandedKey(29) WHEN out0_49 = to_unsigned(16#1E#, 8) ELSE
      expandedKey(30) WHEN out0_49 = to_unsigned(16#1F#, 8) ELSE
      expandedKey(31) WHEN out0_49 = to_unsigned(16#20#, 8) ELSE
      expandedKey(32) WHEN out0_49 = to_unsigned(16#21#, 8) ELSE
      expandedKey(33) WHEN out0_49 = to_unsigned(16#22#, 8) ELSE
      expandedKey(34) WHEN out0_49 = to_unsigned(16#23#, 8) ELSE
      expandedKey(35) WHEN out0_49 = to_unsigned(16#24#, 8) ELSE
      expandedKey(36) WHEN out0_49 = to_unsigned(16#25#, 8) ELSE
      expandedKey(37) WHEN out0_49 = to_unsigned(16#26#, 8) ELSE
      expandedKey(38) WHEN out0_49 = to_unsigned(16#27#, 8) ELSE
      expandedKey(39) WHEN out0_49 = to_unsigned(16#28#, 8) ELSE
      expandedKey(40) WHEN out0_49 = to_unsigned(16#29#, 8) ELSE
      expandedKey(41) WHEN out0_49 = to_unsigned(16#2A#, 8) ELSE
      expandedKey(42) WHEN out0_49 = to_unsigned(16#2B#, 8) ELSE
      expandedKey(43) WHEN out0_49 = to_unsigned(16#2C#, 8) ELSE
      expandedKey(44) WHEN out0_49 = to_unsigned(16#2D#, 8) ELSE
      expandedKey(45) WHEN out0_49 = to_unsigned(16#2E#, 8) ELSE
      expandedKey(46) WHEN out0_49 = to_unsigned(16#2F#, 8) ELSE
      expandedKey(47) WHEN out0_49 = to_unsigned(16#30#, 8) ELSE
      expandedKey(48) WHEN out0_49 = to_unsigned(16#31#, 8) ELSE
      expandedKey(49) WHEN out0_49 = to_unsigned(16#32#, 8) ELSE
      expandedKey(50) WHEN out0_49 = to_unsigned(16#33#, 8) ELSE
      expandedKey(51) WHEN out0_49 = to_unsigned(16#34#, 8) ELSE
      expandedKey(52) WHEN out0_49 = to_unsigned(16#35#, 8) ELSE
      expandedKey(53) WHEN out0_49 = to_unsigned(16#36#, 8) ELSE
      expandedKey(54) WHEN out0_49 = to_unsigned(16#37#, 8) ELSE
      expandedKey(55) WHEN out0_49 = to_unsigned(16#38#, 8) ELSE
      expandedKey(56) WHEN out0_49 = to_unsigned(16#39#, 8) ELSE
      expandedKey(57) WHEN out0_49 = to_unsigned(16#3A#, 8) ELSE
      expandedKey(58) WHEN out0_49 = to_unsigned(16#3B#, 8) ELSE
      expandedKey(59) WHEN out0_49 = to_unsigned(16#3C#, 8) ELSE
      expandedKey(60) WHEN out0_49 = to_unsigned(16#3D#, 8) ELSE
      expandedKey(61) WHEN out0_49 = to_unsigned(16#3E#, 8) ELSE
      expandedKey(62) WHEN out0_49 = to_unsigned(16#3F#, 8) ELSE
      expandedKey(63) WHEN out0_49 = to_unsigned(16#40#, 8) ELSE
      expandedKey(64) WHEN out0_49 = to_unsigned(16#41#, 8) ELSE
      expandedKey(65) WHEN out0_49 = to_unsigned(16#42#, 8) ELSE
      expandedKey(66) WHEN out0_49 = to_unsigned(16#43#, 8) ELSE
      expandedKey(67) WHEN out0_49 = to_unsigned(16#44#, 8) ELSE
      expandedKey(68) WHEN out0_49 = to_unsigned(16#45#, 8) ELSE
      expandedKey(69) WHEN out0_49 = to_unsigned(16#46#, 8) ELSE
      expandedKey(70) WHEN out0_49 = to_unsigned(16#47#, 8) ELSE
      expandedKey(71) WHEN out0_49 = to_unsigned(16#48#, 8) ELSE
      expandedKey(72) WHEN out0_49 = to_unsigned(16#49#, 8) ELSE
      expandedKey(73) WHEN out0_49 = to_unsigned(16#4A#, 8) ELSE
      expandedKey(74) WHEN out0_49 = to_unsigned(16#4B#, 8) ELSE
      expandedKey(75) WHEN out0_49 = to_unsigned(16#4C#, 8) ELSE
      expandedKey(76) WHEN out0_49 = to_unsigned(16#4D#, 8) ELSE
      expandedKey(77) WHEN out0_49 = to_unsigned(16#4E#, 8) ELSE
      expandedKey(78) WHEN out0_49 = to_unsigned(16#4F#, 8) ELSE
      expandedKey(79) WHEN out0_49 = to_unsigned(16#50#, 8) ELSE
      expandedKey(80) WHEN out0_49 = to_unsigned(16#51#, 8) ELSE
      expandedKey(81) WHEN out0_49 = to_unsigned(16#52#, 8) ELSE
      expandedKey(82) WHEN out0_49 = to_unsigned(16#53#, 8) ELSE
      expandedKey(83) WHEN out0_49 = to_unsigned(16#54#, 8) ELSE
      expandedKey(84) WHEN out0_49 = to_unsigned(16#55#, 8) ELSE
      expandedKey(85) WHEN out0_49 = to_unsigned(16#56#, 8) ELSE
      expandedKey(86) WHEN out0_49 = to_unsigned(16#57#, 8) ELSE
      expandedKey(87) WHEN out0_49 = to_unsigned(16#58#, 8) ELSE
      expandedKey(88) WHEN out0_49 = to_unsigned(16#59#, 8) ELSE
      expandedKey(89) WHEN out0_49 = to_unsigned(16#5A#, 8) ELSE
      expandedKey(90) WHEN out0_49 = to_unsigned(16#5B#, 8) ELSE
      expandedKey(91) WHEN out0_49 = to_unsigned(16#5C#, 8) ELSE
      expandedKey(92) WHEN out0_49 = to_unsigned(16#5D#, 8) ELSE
      expandedKey(93) WHEN out0_49 = to_unsigned(16#5E#, 8) ELSE
      expandedKey(94) WHEN out0_49 = to_unsigned(16#5F#, 8) ELSE
      expandedKey(95) WHEN out0_49 = to_unsigned(16#60#, 8) ELSE
      expandedKey(96) WHEN out0_49 = to_unsigned(16#61#, 8) ELSE
      expandedKey(97) WHEN out0_49 = to_unsigned(16#62#, 8) ELSE
      expandedKey(98) WHEN out0_49 = to_unsigned(16#63#, 8) ELSE
      expandedKey(99) WHEN out0_49 = to_unsigned(16#64#, 8) ELSE
      expandedKey(100) WHEN out0_49 = to_unsigned(16#65#, 8) ELSE
      expandedKey(101) WHEN out0_49 = to_unsigned(16#66#, 8) ELSE
      expandedKey(102) WHEN out0_49 = to_unsigned(16#67#, 8) ELSE
      expandedKey(103) WHEN out0_49 = to_unsigned(16#68#, 8) ELSE
      expandedKey(104) WHEN out0_49 = to_unsigned(16#69#, 8) ELSE
      expandedKey(105) WHEN out0_49 = to_unsigned(16#6A#, 8) ELSE
      expandedKey(106) WHEN out0_49 = to_unsigned(16#6B#, 8) ELSE
      expandedKey(107) WHEN out0_49 = to_unsigned(16#6C#, 8) ELSE
      expandedKey(108) WHEN out0_49 = to_unsigned(16#6D#, 8) ELSE
      expandedKey(109) WHEN out0_49 = to_unsigned(16#6E#, 8) ELSE
      expandedKey(110) WHEN out0_49 = to_unsigned(16#6F#, 8) ELSE
      expandedKey(111) WHEN out0_49 = to_unsigned(16#70#, 8) ELSE
      expandedKey(112) WHEN out0_49 = to_unsigned(16#71#, 8) ELSE
      expandedKey(113) WHEN out0_49 = to_unsigned(16#72#, 8) ELSE
      expandedKey(114) WHEN out0_49 = to_unsigned(16#73#, 8) ELSE
      expandedKey(115) WHEN out0_49 = to_unsigned(16#74#, 8) ELSE
      expandedKey(116) WHEN out0_49 = to_unsigned(16#75#, 8) ELSE
      expandedKey(117) WHEN out0_49 = to_unsigned(16#76#, 8) ELSE
      expandedKey(118) WHEN out0_49 = to_unsigned(16#77#, 8) ELSE
      expandedKey(119) WHEN out0_49 = to_unsigned(16#78#, 8) ELSE
      expandedKey(120) WHEN out0_49 = to_unsigned(16#79#, 8) ELSE
      expandedKey(121) WHEN out0_49 = to_unsigned(16#7A#, 8) ELSE
      expandedKey(122) WHEN out0_49 = to_unsigned(16#7B#, 8) ELSE
      expandedKey(123) WHEN out0_49 = to_unsigned(16#7C#, 8) ELSE
      expandedKey(124) WHEN out0_49 = to_unsigned(16#7D#, 8) ELSE
      expandedKey(125) WHEN out0_49 = to_unsigned(16#7E#, 8) ELSE
      expandedKey(126) WHEN out0_49 = to_unsigned(16#7F#, 8) ELSE
      expandedKey(127) WHEN out0_49 = to_unsigned(16#80#, 8) ELSE
      expandedKey(128) WHEN out0_49 = to_unsigned(16#81#, 8) ELSE
      expandedKey(129) WHEN out0_49 = to_unsigned(16#82#, 8) ELSE
      expandedKey(130) WHEN out0_49 = to_unsigned(16#83#, 8) ELSE
      expandedKey(131) WHEN out0_49 = to_unsigned(16#84#, 8) ELSE
      expandedKey(132) WHEN out0_49 = to_unsigned(16#85#, 8) ELSE
      expandedKey(133) WHEN out0_49 = to_unsigned(16#86#, 8) ELSE
      expandedKey(134) WHEN out0_49 = to_unsigned(16#87#, 8) ELSE
      expandedKey(135) WHEN out0_49 = to_unsigned(16#88#, 8) ELSE
      expandedKey(136) WHEN out0_49 = to_unsigned(16#89#, 8) ELSE
      expandedKey(137) WHEN out0_49 = to_unsigned(16#8A#, 8) ELSE
      expandedKey(138) WHEN out0_49 = to_unsigned(16#8B#, 8) ELSE
      expandedKey(139) WHEN out0_49 = to_unsigned(16#8C#, 8) ELSE
      expandedKey(140) WHEN out0_49 = to_unsigned(16#8D#, 8) ELSE
      expandedKey(141) WHEN out0_49 = to_unsigned(16#8E#, 8) ELSE
      expandedKey(142) WHEN out0_49 = to_unsigned(16#8F#, 8) ELSE
      expandedKey(143) WHEN out0_49 = to_unsigned(16#90#, 8) ELSE
      expandedKey(144) WHEN out0_49 = to_unsigned(16#91#, 8) ELSE
      expandedKey(145) WHEN out0_49 = to_unsigned(16#92#, 8) ELSE
      expandedKey(146) WHEN out0_49 = to_unsigned(16#93#, 8) ELSE
      expandedKey(147) WHEN out0_49 = to_unsigned(16#94#, 8) ELSE
      expandedKey(148) WHEN out0_49 = to_unsigned(16#95#, 8) ELSE
      expandedKey(149) WHEN out0_49 = to_unsigned(16#96#, 8) ELSE
      expandedKey(150) WHEN out0_49 = to_unsigned(16#97#, 8) ELSE
      expandedKey(151) WHEN out0_49 = to_unsigned(16#98#, 8) ELSE
      expandedKey(152) WHEN out0_49 = to_unsigned(16#99#, 8) ELSE
      expandedKey(153) WHEN out0_49 = to_unsigned(16#9A#, 8) ELSE
      expandedKey(154) WHEN out0_49 = to_unsigned(16#9B#, 8) ELSE
      expandedKey(155) WHEN out0_49 = to_unsigned(16#9C#, 8) ELSE
      expandedKey(156) WHEN out0_49 = to_unsigned(16#9D#, 8) ELSE
      expandedKey(157) WHEN out0_49 = to_unsigned(16#9E#, 8) ELSE
      expandedKey(158) WHEN out0_49 = to_unsigned(16#9F#, 8) ELSE
      expandedKey(159) WHEN out0_49 = to_unsigned(16#A0#, 8) ELSE
      expandedKey(160) WHEN out0_49 = to_unsigned(16#A1#, 8) ELSE
      expandedKey(161) WHEN out0_49 = to_unsigned(16#A2#, 8) ELSE
      expandedKey(162) WHEN out0_49 = to_unsigned(16#A3#, 8) ELSE
      expandedKey(163) WHEN out0_49 = to_unsigned(16#A4#, 8) ELSE
      expandedKey(164) WHEN out0_49 = to_unsigned(16#A5#, 8) ELSE
      expandedKey(165) WHEN out0_49 = to_unsigned(16#A6#, 8) ELSE
      expandedKey(166) WHEN out0_49 = to_unsigned(16#A7#, 8) ELSE
      expandedKey(167) WHEN out0_49 = to_unsigned(16#A8#, 8) ELSE
      expandedKey(168) WHEN out0_49 = to_unsigned(16#A9#, 8) ELSE
      expandedKey(169) WHEN out0_49 = to_unsigned(16#AA#, 8) ELSE
      expandedKey(170) WHEN out0_49 = to_unsigned(16#AB#, 8) ELSE
      expandedKey(171) WHEN out0_49 = to_unsigned(16#AC#, 8) ELSE
      expandedKey(172) WHEN out0_49 = to_unsigned(16#AD#, 8) ELSE
      expandedKey(173) WHEN out0_49 = to_unsigned(16#AE#, 8) ELSE
      expandedKey(174) WHEN out0_49 = to_unsigned(16#AF#, 8) ELSE
      expandedKey(175) WHEN out0_49 = to_unsigned(16#B0#, 8) ELSE
      expandedKey(176) WHEN out0_49 = to_unsigned(16#B1#, 8) ELSE
      expandedKey(177) WHEN out0_49 = to_unsigned(16#B2#, 8) ELSE
      expandedKey(178) WHEN out0_49 = to_unsigned(16#B3#, 8) ELSE
      expandedKey(179) WHEN out0_49 = to_unsigned(16#B4#, 8) ELSE
      expandedKey(180) WHEN out0_49 = to_unsigned(16#B5#, 8) ELSE
      expandedKey(181) WHEN out0_49 = to_unsigned(16#B6#, 8) ELSE
      expandedKey(182) WHEN out0_49 = to_unsigned(16#B7#, 8) ELSE
      expandedKey(183) WHEN out0_49 = to_unsigned(16#B8#, 8) ELSE
      expandedKey(184) WHEN out0_49 = to_unsigned(16#B9#, 8) ELSE
      expandedKey(185) WHEN out0_49 = to_unsigned(16#BA#, 8) ELSE
      expandedKey(186) WHEN out0_49 = to_unsigned(16#BB#, 8) ELSE
      expandedKey(187) WHEN out0_49 = to_unsigned(16#BC#, 8) ELSE
      expandedKey(188) WHEN out0_49 = to_unsigned(16#BD#, 8) ELSE
      expandedKey(189) WHEN out0_49 = to_unsigned(16#BE#, 8) ELSE
      expandedKey(190) WHEN out0_49 = to_unsigned(16#BF#, 8) ELSE
      expandedKey(191) WHEN out0_49 = to_unsigned(16#C0#, 8) ELSE
      expandedKey(192) WHEN out0_49 = to_unsigned(16#C1#, 8) ELSE
      expandedKey(193) WHEN out0_49 = to_unsigned(16#C2#, 8) ELSE
      expandedKey(194) WHEN out0_49 = to_unsigned(16#C3#, 8) ELSE
      expandedKey(195) WHEN out0_49 = to_unsigned(16#C4#, 8) ELSE
      expandedKey(196) WHEN out0_49 = to_unsigned(16#C5#, 8) ELSE
      expandedKey(197) WHEN out0_49 = to_unsigned(16#C6#, 8) ELSE
      expandedKey(198) WHEN out0_49 = to_unsigned(16#C7#, 8) ELSE
      expandedKey(199) WHEN out0_49 = to_unsigned(16#C8#, 8) ELSE
      expandedKey(200) WHEN out0_49 = to_unsigned(16#C9#, 8) ELSE
      expandedKey(201) WHEN out0_49 = to_unsigned(16#CA#, 8) ELSE
      expandedKey(202) WHEN out0_49 = to_unsigned(16#CB#, 8) ELSE
      expandedKey(203) WHEN out0_49 = to_unsigned(16#CC#, 8) ELSE
      expandedKey(204) WHEN out0_49 = to_unsigned(16#CD#, 8) ELSE
      expandedKey(205) WHEN out0_49 = to_unsigned(16#CE#, 8) ELSE
      expandedKey(206) WHEN out0_49 = to_unsigned(16#CF#, 8) ELSE
      expandedKey(207) WHEN out0_49 = to_unsigned(16#D0#, 8) ELSE
      expandedKey(208) WHEN out0_49 = to_unsigned(16#D1#, 8) ELSE
      expandedKey(209) WHEN out0_49 = to_unsigned(16#D2#, 8) ELSE
      expandedKey(210) WHEN out0_49 = to_unsigned(16#D3#, 8) ELSE
      expandedKey(211) WHEN out0_49 = to_unsigned(16#D4#, 8) ELSE
      expandedKey(212) WHEN out0_49 = to_unsigned(16#D5#, 8) ELSE
      expandedKey(213) WHEN out0_49 = to_unsigned(16#D6#, 8) ELSE
      expandedKey(214) WHEN out0_49 = to_unsigned(16#D7#, 8) ELSE
      expandedKey(215) WHEN out0_49 = to_unsigned(16#D8#, 8) ELSE
      expandedKey(216) WHEN out0_49 = to_unsigned(16#D9#, 8) ELSE
      expandedKey(217) WHEN out0_49 = to_unsigned(16#DA#, 8) ELSE
      expandedKey(218) WHEN out0_49 = to_unsigned(16#DB#, 8) ELSE
      expandedKey(219) WHEN out0_49 = to_unsigned(16#DC#, 8) ELSE
      expandedKey(220) WHEN out0_49 = to_unsigned(16#DD#, 8) ELSE
      expandedKey(221) WHEN out0_49 = to_unsigned(16#DE#, 8) ELSE
      expandedKey(222) WHEN out0_49 = to_unsigned(16#DF#, 8) ELSE
      expandedKey(223) WHEN out0_49 = to_unsigned(16#E0#, 8) ELSE
      expandedKey(224) WHEN out0_49 = to_unsigned(16#E1#, 8) ELSE
      expandedKey(225) WHEN out0_49 = to_unsigned(16#E2#, 8) ELSE
      expandedKey(226) WHEN out0_49 = to_unsigned(16#E3#, 8) ELSE
      expandedKey(227) WHEN out0_49 = to_unsigned(16#E4#, 8) ELSE
      expandedKey(228) WHEN out0_49 = to_unsigned(16#E5#, 8) ELSE
      expandedKey(229) WHEN out0_49 = to_unsigned(16#E6#, 8) ELSE
      expandedKey(230) WHEN out0_49 = to_unsigned(16#E7#, 8) ELSE
      expandedKey(231) WHEN out0_49 = to_unsigned(16#E8#, 8) ELSE
      expandedKey(232) WHEN out0_49 = to_unsigned(16#E9#, 8) ELSE
      expandedKey(233) WHEN out0_49 = to_unsigned(16#EA#, 8) ELSE
      expandedKey(234) WHEN out0_49 = to_unsigned(16#EB#, 8) ELSE
      expandedKey(235) WHEN out0_49 = to_unsigned(16#EC#, 8) ELSE
      expandedKey(236) WHEN out0_49 = to_unsigned(16#ED#, 8) ELSE
      expandedKey(237) WHEN out0_49 = to_unsigned(16#EE#, 8) ELSE
      expandedKey(238) WHEN out0_49 = to_unsigned(16#EF#, 8) ELSE
      expandedKey(239);

  
  out0_114(0) <= ss(0) WHEN out0_10 = '0' ELSE
      ss(0);
  
  out0_114(1) <= ss(1) WHEN out0_10 = '0' ELSE
      ss(1);
  
  out0_114(2) <= ss(2) WHEN out0_10 = '0' ELSE
      ss(2);
  
  out0_114(3) <= ss(3) WHEN out0_10 = '0' ELSE
      ss(3);
  
  out0_114(4) <= ss(4) WHEN out0_10 = '0' ELSE
      ss(4);
  
  out0_114(5) <= ss(5) WHEN out0_10 = '0' ELSE
      ss(5);
  
  out0_114(6) <= ss(6) WHEN out0_10 = '0' ELSE
      ss(6);
  
  out0_114(7) <= ss(7) WHEN out0_10 = '0' ELSE
      ss(7);
  
  out0_114(8) <= ss(8) WHEN out0_10 = '0' ELSE
      ss(8);
  
  out0_114(9) <= ss(9) WHEN out0_10 = '0' ELSE
      ss(9);
  
  out0_114(10) <= ss(10) WHEN out0_10 = '0' ELSE
      ss(10);
  
  out0_114(11) <= ss(11) WHEN out0_10 = '0' ELSE
      ss(11);
  
  out0_114(12) <= ss(12) WHEN out0_10 = '0' ELSE
      ss(12);
  
  out0_114(13) <= ss(13) WHEN out0_10 = '0' ELSE
      ss(13);
  
  out0_114(14) <= ss(14) WHEN out0_10 = '0' ELSE
      ss(14);
  
  out0_114(15) <= ss(15) WHEN out0_10 = '0' ELSE
      ss(15);

  
  out0_115(0) <= out0_114(0) WHEN out0_12 = '0' ELSE
      ss_1(0);
  
  out0_115(1) <= out0_114(1) WHEN out0_12 = '0' ELSE
      ss_1(1);
  
  out0_115(2) <= out0_114(2) WHEN out0_12 = '0' ELSE
      ss_1(2);
  
  out0_115(3) <= out0_114(3) WHEN out0_12 = '0' ELSE
      ss_1(3);
  
  out0_115(4) <= out0_114(4) WHEN out0_12 = '0' ELSE
      ss_1(4);
  
  out0_115(5) <= out0_114(5) WHEN out0_12 = '0' ELSE
      ss_1(5);
  
  out0_115(6) <= out0_114(6) WHEN out0_12 = '0' ELSE
      ss_1(6);
  
  out0_115(7) <= out0_114(7) WHEN out0_12 = '0' ELSE
      ss_1(7);
  
  out0_115(8) <= out0_114(8) WHEN out0_12 = '0' ELSE
      ss_1(8);
  
  out0_115(9) <= out0_114(9) WHEN out0_12 = '0' ELSE
      ss_1(9);
  
  out0_115(10) <= out0_114(10) WHEN out0_12 = '0' ELSE
      ss_1(10);
  
  out0_115(11) <= out0_114(11) WHEN out0_12 = '0' ELSE
      ss_1(11);
  
  out0_115(12) <= out0_114(12) WHEN out0_12 = '0' ELSE
      ss_1(12);
  
  out0_115(13) <= out0_114(13) WHEN out0_12 = '0' ELSE
      ss_1(13);
  
  out0_115(14) <= out0_114(14) WHEN out0_12 = '0' ELSE
      ss_1(14);
  
  out0_115(15) <= out0_114(15) WHEN out0_12 = '0' ELSE
      ss_1(15);

  
  out0_116(0) <= out0_115(0) WHEN out0_14 = '0' ELSE
      ss(0);
  
  out0_116(1) <= out0_115(1) WHEN out0_14 = '0' ELSE
      ss(1);
  
  out0_116(2) <= out0_115(2) WHEN out0_14 = '0' ELSE
      ss(2);
  
  out0_116(3) <= out0_115(3) WHEN out0_14 = '0' ELSE
      ss(3);
  
  out0_116(4) <= out0_115(4) WHEN out0_14 = '0' ELSE
      ss(4);
  
  out0_116(5) <= out0_115(5) WHEN out0_14 = '0' ELSE
      ss(5);
  
  out0_116(6) <= out0_115(6) WHEN out0_14 = '0' ELSE
      ss(6);
  
  out0_116(7) <= out0_115(7) WHEN out0_14 = '0' ELSE
      ss(7);
  
  out0_116(8) <= out0_115(8) WHEN out0_14 = '0' ELSE
      ss(8);
  
  out0_116(9) <= out0_115(9) WHEN out0_14 = '0' ELSE
      ss(9);
  
  out0_116(10) <= out0_115(10) WHEN out0_14 = '0' ELSE
      ss(10);
  
  out0_116(11) <= out0_115(11) WHEN out0_14 = '0' ELSE
      ss(11);
  
  out0_116(12) <= out0_115(12) WHEN out0_14 = '0' ELSE
      ss(12);
  
  out0_116(13) <= out0_115(13) WHEN out0_14 = '0' ELSE
      ss(13);
  
  out0_116(14) <= out0_115(14) WHEN out0_14 = '0' ELSE
      ss(14);
  
  out0_116(15) <= out0_115(15) WHEN out0_14 = '0' ELSE
      ss(15);

  
  out0_117(0) <= out0_116(0) WHEN out0_16 = '0' ELSE
      ss(0);
  
  out0_117(1) <= out0_116(1) WHEN out0_16 = '0' ELSE
      ss(1);
  
  out0_117(2) <= out0_116(2) WHEN out0_16 = '0' ELSE
      ss(2);
  
  out0_117(3) <= out0_116(3) WHEN out0_16 = '0' ELSE
      ss(3);
  
  out0_117(4) <= out0_116(4) WHEN out0_16 = '0' ELSE
      ss(4);
  
  out0_117(5) <= out0_116(5) WHEN out0_16 = '0' ELSE
      ss(5);
  
  out0_117(6) <= out0_116(6) WHEN out0_16 = '0' ELSE
      ss(6);
  
  out0_117(7) <= out0_116(7) WHEN out0_16 = '0' ELSE
      ss(7);
  
  out0_117(8) <= out0_116(8) WHEN out0_16 = '0' ELSE
      ss(8);
  
  out0_117(9) <= out0_116(9) WHEN out0_16 = '0' ELSE
      ss(9);
  
  out0_117(10) <= out0_116(10) WHEN out0_16 = '0' ELSE
      ss(10);
  
  out0_117(11) <= out0_116(11) WHEN out0_16 = '0' ELSE
      ss(11);
  
  out0_117(12) <= out0_116(12) WHEN out0_16 = '0' ELSE
      ss(12);
  
  out0_117(13) <= out0_116(13) WHEN out0_16 = '0' ELSE
      ss(13);
  
  out0_117(14) <= out0_116(14) WHEN out0_16 = '0' ELSE
      ss(14);
  
  out0_117(15) <= out0_116(15) WHEN out0_16 = '0' ELSE
      ss(15);

  
  out0_118(0) <= out0_117(0) WHEN out0_18 = '0' ELSE
      ss(0);
  
  out0_118(1) <= out0_117(1) WHEN out0_18 = '0' ELSE
      ss(1);
  
  out0_118(2) <= out0_117(2) WHEN out0_18 = '0' ELSE
      ss(2);
  
  out0_118(3) <= out0_117(3) WHEN out0_18 = '0' ELSE
      ss(3);
  
  out0_118(4) <= out0_117(4) WHEN out0_18 = '0' ELSE
      ss(4);
  
  out0_118(5) <= out0_117(5) WHEN out0_18 = '0' ELSE
      ss(5);
  
  out0_118(6) <= out0_117(6) WHEN out0_18 = '0' ELSE
      ss(6);
  
  out0_118(7) <= out0_117(7) WHEN out0_18 = '0' ELSE
      ss(7);
  
  out0_118(8) <= out0_117(8) WHEN out0_18 = '0' ELSE
      ss(8);
  
  out0_118(9) <= out0_117(9) WHEN out0_18 = '0' ELSE
      ss(9);
  
  out0_118(10) <= out0_117(10) WHEN out0_18 = '0' ELSE
      ss(10);
  
  out0_118(11) <= out0_117(11) WHEN out0_18 = '0' ELSE
      ss(11);
  
  out0_118(12) <= out0_117(12) WHEN out0_18 = '0' ELSE
      ss(12);
  
  out0_118(13) <= out0_117(13) WHEN out0_18 = '0' ELSE
      ss(13);
  
  out0_118(14) <= out0_117(14) WHEN out0_18 = '0' ELSE
      ss(14);
  
  out0_118(15) <= out0_117(15) WHEN out0_18 = '0' ELSE
      ss(15);

  
  out0_119(0) <= out0_118(0) WHEN out0_20 = '0' ELSE
      ss(0);
  
  out0_119(1) <= out0_118(1) WHEN out0_20 = '0' ELSE
      ss(1);
  
  out0_119(2) <= out0_118(2) WHEN out0_20 = '0' ELSE
      ss(2);
  
  out0_119(3) <= out0_118(3) WHEN out0_20 = '0' ELSE
      ss(3);
  
  out0_119(4) <= out0_118(4) WHEN out0_20 = '0' ELSE
      ss(4);
  
  out0_119(5) <= out0_118(5) WHEN out0_20 = '0' ELSE
      ss(5);
  
  out0_119(6) <= out0_118(6) WHEN out0_20 = '0' ELSE
      ss(6);
  
  out0_119(7) <= out0_118(7) WHEN out0_20 = '0' ELSE
      ss(7);
  
  out0_119(8) <= out0_118(8) WHEN out0_20 = '0' ELSE
      ss(8);
  
  out0_119(9) <= out0_118(9) WHEN out0_20 = '0' ELSE
      ss(9);
  
  out0_119(10) <= out0_118(10) WHEN out0_20 = '0' ELSE
      ss(10);
  
  out0_119(11) <= out0_118(11) WHEN out0_20 = '0' ELSE
      ss(11);
  
  out0_119(12) <= out0_118(12) WHEN out0_20 = '0' ELSE
      ss(12);
  
  out0_119(13) <= out0_118(13) WHEN out0_20 = '0' ELSE
      ss(13);
  
  out0_119(14) <= out0_118(14) WHEN out0_20 = '0' ELSE
      ss(14);
  
  out0_119(15) <= out0_118(15) WHEN out0_20 = '0' ELSE
      ss(15);

  
  out0_120(0) <= out0_119(0) WHEN out0_22 = '0' ELSE
      ss(0);
  
  out0_120(1) <= out0_119(1) WHEN out0_22 = '0' ELSE
      ss(1);
  
  out0_120(2) <= out0_119(2) WHEN out0_22 = '0' ELSE
      ss(2);
  
  out0_120(3) <= out0_119(3) WHEN out0_22 = '0' ELSE
      ss(3);
  
  out0_120(4) <= out0_119(4) WHEN out0_22 = '0' ELSE
      ss(4);
  
  out0_120(5) <= out0_119(5) WHEN out0_22 = '0' ELSE
      ss(5);
  
  out0_120(6) <= out0_119(6) WHEN out0_22 = '0' ELSE
      ss(6);
  
  out0_120(7) <= out0_119(7) WHEN out0_22 = '0' ELSE
      ss(7);
  
  out0_120(8) <= out0_119(8) WHEN out0_22 = '0' ELSE
      ss(8);
  
  out0_120(9) <= out0_119(9) WHEN out0_22 = '0' ELSE
      ss(9);
  
  out0_120(10) <= out0_119(10) WHEN out0_22 = '0' ELSE
      ss(10);
  
  out0_120(11) <= out0_119(11) WHEN out0_22 = '0' ELSE
      ss(11);
  
  out0_120(12) <= out0_119(12) WHEN out0_22 = '0' ELSE
      ss(12);
  
  out0_120(13) <= out0_119(13) WHEN out0_22 = '0' ELSE
      ss(13);
  
  out0_120(14) <= out0_119(14) WHEN out0_22 = '0' ELSE
      ss(14);
  
  out0_120(15) <= out0_119(15) WHEN out0_22 = '0' ELSE
      ss(15);

  
  ss_2(0) <= out0_120(0) WHEN out0_24 = '0' ELSE
      ss(0);
  
  ss_2(1) <= out0_120(1) WHEN out0_24 = '0' ELSE
      ss(1);
  
  ss_2(2) <= out0_120(2) WHEN out0_24 = '0' ELSE
      ss(2);
  
  ss_2(3) <= out0_120(3) WHEN out0_24 = '0' ELSE
      ss(3);
  
  ss_2(4) <= out0_120(4) WHEN out0_24 = '0' ELSE
      ss(4);
  
  ss_2(5) <= out0_120(5) WHEN out0_24 = '0' ELSE
      ss(5);
  
  ss_2(6) <= out0_120(6) WHEN out0_24 = '0' ELSE
      ss(6);
  
  ss_2(7) <= out0_120(7) WHEN out0_24 = '0' ELSE
      ss(7);
  
  ss_2(8) <= out0_120(8) WHEN out0_24 = '0' ELSE
      ss(8);
  
  ss_2(9) <= out0_120(9) WHEN out0_24 = '0' ELSE
      ss(9);
  
  ss_2(10) <= out0_120(10) WHEN out0_24 = '0' ELSE
      ss(10);
  
  ss_2(11) <= out0_120(11) WHEN out0_24 = '0' ELSE
      ss(11);
  
  ss_2(12) <= out0_120(12) WHEN out0_24 = '0' ELSE
      ss(12);
  
  ss_2(13) <= out0_120(13) WHEN out0_24 = '0' ELSE
      ss(13);
  
  ss_2(14) <= out0_120(14) WHEN out0_24 = '0' ELSE
      ss(14);
  
  ss_2(15) <= out0_120(15) WHEN out0_24 = '0' ELSE
      ss(15);

  intdelay4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        ss(0) <= to_unsigned(16#00#, 8);
        ss(1) <= to_unsigned(16#00#, 8);
        ss(2) <= to_unsigned(16#00#, 8);
        ss(3) <= to_unsigned(16#00#, 8);
        ss(4) <= to_unsigned(16#00#, 8);
        ss(5) <= to_unsigned(16#00#, 8);
        ss(6) <= to_unsigned(16#00#, 8);
        ss(7) <= to_unsigned(16#00#, 8);
        ss(8) <= to_unsigned(16#00#, 8);
        ss(9) <= to_unsigned(16#00#, 8);
        ss(10) <= to_unsigned(16#00#, 8);
        ss(11) <= to_unsigned(16#00#, 8);
        ss(12) <= to_unsigned(16#00#, 8);
        ss(13) <= to_unsigned(16#00#, 8);
        ss(14) <= to_unsigned(16#00#, 8);
        ss(15) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        ss(0) <= ss_2(0);
        ss(1) <= ss_2(1);
        ss(2) <= ss_2(2);
        ss(3) <= ss_2(3);
        ss(4) <= ss_2(4);
        ss(5) <= ss_2(5);
        ss(6) <= ss_2(6);
        ss(7) <= ss_2(7);
        ss(8) <= ss_2(8);
        ss(9) <= ss_2(9);
        ss(10) <= ss_2(10);
        ss(11) <= ss_2(11);
        ss(12) <= ss_2(12);
        ss(13) <= ss_2(13);
        ss(14) <= ss_2(14);
        ss(15) <= ss_2(15);
      END IF;
    END IF;
  END PROCESS intdelay4_process;


  
  ss_1(0) <= out0_113 WHEN ii_8 = to_unsigned(16#01#, 8) ELSE
      ss(0);
  
  ss_1(1) <= out0_113 WHEN ii_8 = to_unsigned(16#02#, 8) ELSE
      ss(1);
  
  ss_1(2) <= out0_113 WHEN ii_8 = to_unsigned(16#03#, 8) ELSE
      ss(2);
  
  ss_1(3) <= out0_113 WHEN ii_8 = to_unsigned(16#04#, 8) ELSE
      ss(3);
  
  ss_1(4) <= out0_113 WHEN ii_8 = to_unsigned(16#05#, 8) ELSE
      ss(4);
  
  ss_1(5) <= out0_113 WHEN ii_8 = to_unsigned(16#06#, 8) ELSE
      ss(5);
  
  ss_1(6) <= out0_113 WHEN ii_8 = to_unsigned(16#07#, 8) ELSE
      ss(6);
  
  ss_1(7) <= out0_113 WHEN ii_8 = to_unsigned(16#08#, 8) ELSE
      ss(7);
  
  ss_1(8) <= out0_113 WHEN ii_8 = to_unsigned(16#09#, 8) ELSE
      ss(8);
  
  ss_1(9) <= out0_113 WHEN ii_8 = to_unsigned(16#0A#, 8) ELSE
      ss(9);
  
  ss_1(10) <= out0_113 WHEN ii_8 = to_unsigned(16#0B#, 8) ELSE
      ss(10);
  
  ss_1(11) <= out0_113 WHEN ii_8 = to_unsigned(16#0C#, 8) ELSE
      ss(11);
  
  ss_1(12) <= out0_113 WHEN ii_8 = to_unsigned(16#0D#, 8) ELSE
      ss(12);
  
  ss_1(13) <= out0_113 WHEN ii_8 = to_unsigned(16#0E#, 8) ELSE
      ss(13);
  
  ss_1(14) <= out0_113 WHEN ii_8 = to_unsigned(16#0F#, 8) ELSE
      ss(14);
  
  ss_1(15) <= out0_113 WHEN ii_8 = to_unsigned(16#10#, 8) ELSE
      ss(15);

  
  out0_121 <= ss_1(0) WHEN ii_8 = to_unsigned(16#01#, 8) ELSE
      ss_1(1) WHEN ii_8 = to_unsigned(16#02#, 8) ELSE
      ss_1(2) WHEN ii_8 = to_unsigned(16#03#, 8) ELSE
      ss_1(3) WHEN ii_8 = to_unsigned(16#04#, 8) ELSE
      ss_1(4) WHEN ii_8 = to_unsigned(16#05#, 8) ELSE
      ss_1(5) WHEN ii_8 = to_unsigned(16#06#, 8) ELSE
      ss_1(6) WHEN ii_8 = to_unsigned(16#07#, 8) ELSE
      ss_1(7) WHEN ii_8 = to_unsigned(16#08#, 8) ELSE
      ss_1(8) WHEN ii_8 = to_unsigned(16#09#, 8) ELSE
      ss_1(9) WHEN ii_8 = to_unsigned(16#0A#, 8) ELSE
      ss_1(10) WHEN ii_8 = to_unsigned(16#0B#, 8) ELSE
      ss_1(11) WHEN ii_8 = to_unsigned(16#0C#, 8) ELSE
      ss_1(12) WHEN ii_8 = to_unsigned(16#0D#, 8) ELSE
      ss_1(13) WHEN ii_8 = to_unsigned(16#0E#, 8) ELSE
      ss_1(14) WHEN ii_8 = to_unsigned(16#0F#, 8) ELSE
      ss_1(15);

  gmul2(0) <= to_unsigned(16#02#, 8);
  gmul2(1) <= to_unsigned(16#04#, 8);
  gmul2(2) <= to_unsigned(16#06#, 8);
  gmul2(3) <= to_unsigned(16#08#, 8);
  gmul2(4) <= to_unsigned(16#0A#, 8);
  gmul2(5) <= to_unsigned(16#0C#, 8);
  gmul2(6) <= to_unsigned(16#0E#, 8);
  gmul2(7) <= to_unsigned(16#10#, 8);
  gmul2(8) <= to_unsigned(16#12#, 8);
  gmul2(9) <= to_unsigned(16#14#, 8);
  gmul2(10) <= to_unsigned(16#16#, 8);
  gmul2(11) <= to_unsigned(16#18#, 8);
  gmul2(12) <= to_unsigned(16#1A#, 8);
  gmul2(13) <= to_unsigned(16#1C#, 8);
  gmul2(14) <= to_unsigned(16#1E#, 8);
  gmul2(15) <= to_unsigned(16#20#, 8);
  gmul2(16) <= to_unsigned(16#22#, 8);
  gmul2(17) <= to_unsigned(16#24#, 8);
  gmul2(18) <= to_unsigned(16#26#, 8);
  gmul2(19) <= to_unsigned(16#28#, 8);
  gmul2(20) <= to_unsigned(16#2A#, 8);
  gmul2(21) <= to_unsigned(16#2C#, 8);
  gmul2(22) <= to_unsigned(16#2E#, 8);
  gmul2(23) <= to_unsigned(16#30#, 8);
  gmul2(24) <= to_unsigned(16#32#, 8);
  gmul2(25) <= to_unsigned(16#34#, 8);
  gmul2(26) <= to_unsigned(16#36#, 8);
  gmul2(27) <= to_unsigned(16#38#, 8);
  gmul2(28) <= to_unsigned(16#3A#, 8);
  gmul2(29) <= to_unsigned(16#3C#, 8);
  gmul2(30) <= to_unsigned(16#3E#, 8);
  gmul2(31) <= to_unsigned(16#40#, 8);
  gmul2(32) <= to_unsigned(16#42#, 8);
  gmul2(33) <= to_unsigned(16#44#, 8);
  gmul2(34) <= to_unsigned(16#46#, 8);
  gmul2(35) <= to_unsigned(16#48#, 8);
  gmul2(36) <= to_unsigned(16#4A#, 8);
  gmul2(37) <= to_unsigned(16#4C#, 8);
  gmul2(38) <= to_unsigned(16#4E#, 8);
  gmul2(39) <= to_unsigned(16#50#, 8);
  gmul2(40) <= to_unsigned(16#52#, 8);
  gmul2(41) <= to_unsigned(16#54#, 8);
  gmul2(42) <= to_unsigned(16#56#, 8);
  gmul2(43) <= to_unsigned(16#58#, 8);
  gmul2(44) <= to_unsigned(16#5A#, 8);
  gmul2(45) <= to_unsigned(16#5C#, 8);
  gmul2(46) <= to_unsigned(16#5E#, 8);
  gmul2(47) <= to_unsigned(16#60#, 8);
  gmul2(48) <= to_unsigned(16#62#, 8);
  gmul2(49) <= to_unsigned(16#64#, 8);
  gmul2(50) <= to_unsigned(16#66#, 8);
  gmul2(51) <= to_unsigned(16#68#, 8);
  gmul2(52) <= to_unsigned(16#6A#, 8);
  gmul2(53) <= to_unsigned(16#6C#, 8);
  gmul2(54) <= to_unsigned(16#6E#, 8);
  gmul2(55) <= to_unsigned(16#70#, 8);
  gmul2(56) <= to_unsigned(16#72#, 8);
  gmul2(57) <= to_unsigned(16#74#, 8);
  gmul2(58) <= to_unsigned(16#76#, 8);
  gmul2(59) <= to_unsigned(16#78#, 8);
  gmul2(60) <= to_unsigned(16#7A#, 8);
  gmul2(61) <= to_unsigned(16#7C#, 8);
  gmul2(62) <= to_unsigned(16#7E#, 8);
  gmul2(63) <= to_unsigned(16#80#, 8);
  gmul2(64) <= to_unsigned(16#82#, 8);
  gmul2(65) <= to_unsigned(16#84#, 8);
  gmul2(66) <= to_unsigned(16#86#, 8);
  gmul2(67) <= to_unsigned(16#88#, 8);
  gmul2(68) <= to_unsigned(16#8A#, 8);
  gmul2(69) <= to_unsigned(16#8C#, 8);
  gmul2(70) <= to_unsigned(16#8E#, 8);
  gmul2(71) <= to_unsigned(16#90#, 8);
  gmul2(72) <= to_unsigned(16#92#, 8);
  gmul2(73) <= to_unsigned(16#94#, 8);
  gmul2(74) <= to_unsigned(16#96#, 8);
  gmul2(75) <= to_unsigned(16#98#, 8);
  gmul2(76) <= to_unsigned(16#9A#, 8);
  gmul2(77) <= to_unsigned(16#9C#, 8);
  gmul2(78) <= to_unsigned(16#9E#, 8);
  gmul2(79) <= to_unsigned(16#A0#, 8);
  gmul2(80) <= to_unsigned(16#A2#, 8);
  gmul2(81) <= to_unsigned(16#A4#, 8);
  gmul2(82) <= to_unsigned(16#A6#, 8);
  gmul2(83) <= to_unsigned(16#A8#, 8);
  gmul2(84) <= to_unsigned(16#AA#, 8);
  gmul2(85) <= to_unsigned(16#AC#, 8);
  gmul2(86) <= to_unsigned(16#AE#, 8);
  gmul2(87) <= to_unsigned(16#B0#, 8);
  gmul2(88) <= to_unsigned(16#B2#, 8);
  gmul2(89) <= to_unsigned(16#B4#, 8);
  gmul2(90) <= to_unsigned(16#B6#, 8);
  gmul2(91) <= to_unsigned(16#B8#, 8);
  gmul2(92) <= to_unsigned(16#BA#, 8);
  gmul2(93) <= to_unsigned(16#BC#, 8);
  gmul2(94) <= to_unsigned(16#BE#, 8);
  gmul2(95) <= to_unsigned(16#C0#, 8);
  gmul2(96) <= to_unsigned(16#C2#, 8);
  gmul2(97) <= to_unsigned(16#C4#, 8);
  gmul2(98) <= to_unsigned(16#C6#, 8);
  gmul2(99) <= to_unsigned(16#C8#, 8);
  gmul2(100) <= to_unsigned(16#CA#, 8);
  gmul2(101) <= to_unsigned(16#CC#, 8);
  gmul2(102) <= to_unsigned(16#CE#, 8);
  gmul2(103) <= to_unsigned(16#D0#, 8);
  gmul2(104) <= to_unsigned(16#D2#, 8);
  gmul2(105) <= to_unsigned(16#D4#, 8);
  gmul2(106) <= to_unsigned(16#D6#, 8);
  gmul2(107) <= to_unsigned(16#D8#, 8);
  gmul2(108) <= to_unsigned(16#DA#, 8);
  gmul2(109) <= to_unsigned(16#DC#, 8);
  gmul2(110) <= to_unsigned(16#DE#, 8);
  gmul2(111) <= to_unsigned(16#E0#, 8);
  gmul2(112) <= to_unsigned(16#E2#, 8);
  gmul2(113) <= to_unsigned(16#E4#, 8);
  gmul2(114) <= to_unsigned(16#E6#, 8);
  gmul2(115) <= to_unsigned(16#E8#, 8);
  gmul2(116) <= to_unsigned(16#EA#, 8);
  gmul2(117) <= to_unsigned(16#EC#, 8);
  gmul2(118) <= to_unsigned(16#EE#, 8);
  gmul2(119) <= to_unsigned(16#F0#, 8);
  gmul2(120) <= to_unsigned(16#F2#, 8);
  gmul2(121) <= to_unsigned(16#F4#, 8);
  gmul2(122) <= to_unsigned(16#F6#, 8);
  gmul2(123) <= to_unsigned(16#F8#, 8);
  gmul2(124) <= to_unsigned(16#FA#, 8);
  gmul2(125) <= to_unsigned(16#FC#, 8);
  gmul2(126) <= to_unsigned(16#FE#, 8);
  gmul2(127) <= to_unsigned(16#1B#, 8);
  gmul2(128) <= to_unsigned(16#19#, 8);
  gmul2(129) <= to_unsigned(16#1F#, 8);
  gmul2(130) <= to_unsigned(16#1D#, 8);
  gmul2(131) <= to_unsigned(16#13#, 8);
  gmul2(132) <= to_unsigned(16#11#, 8);
  gmul2(133) <= to_unsigned(16#17#, 8);
  gmul2(134) <= to_unsigned(16#15#, 8);
  gmul2(135) <= to_unsigned(16#0B#, 8);
  gmul2(136) <= to_unsigned(16#09#, 8);
  gmul2(137) <= to_unsigned(16#0F#, 8);
  gmul2(138) <= to_unsigned(16#0D#, 8);
  gmul2(139) <= to_unsigned(16#03#, 8);
  gmul2(140) <= to_unsigned(16#01#, 8);
  gmul2(141) <= to_unsigned(16#07#, 8);
  gmul2(142) <= to_unsigned(16#05#, 8);
  gmul2(143) <= to_unsigned(16#3B#, 8);
  gmul2(144) <= to_unsigned(16#39#, 8);
  gmul2(145) <= to_unsigned(16#3F#, 8);
  gmul2(146) <= to_unsigned(16#3D#, 8);
  gmul2(147) <= to_unsigned(16#33#, 8);
  gmul2(148) <= to_unsigned(16#31#, 8);
  gmul2(149) <= to_unsigned(16#37#, 8);
  gmul2(150) <= to_unsigned(16#35#, 8);
  gmul2(151) <= to_unsigned(16#2B#, 8);
  gmul2(152) <= to_unsigned(16#29#, 8);
  gmul2(153) <= to_unsigned(16#2F#, 8);
  gmul2(154) <= to_unsigned(16#2D#, 8);
  gmul2(155) <= to_unsigned(16#23#, 8);
  gmul2(156) <= to_unsigned(16#21#, 8);
  gmul2(157) <= to_unsigned(16#27#, 8);
  gmul2(158) <= to_unsigned(16#25#, 8);
  gmul2(159) <= to_unsigned(16#5B#, 8);
  gmul2(160) <= to_unsigned(16#59#, 8);
  gmul2(161) <= to_unsigned(16#5F#, 8);
  gmul2(162) <= to_unsigned(16#5D#, 8);
  gmul2(163) <= to_unsigned(16#53#, 8);
  gmul2(164) <= to_unsigned(16#51#, 8);
  gmul2(165) <= to_unsigned(16#57#, 8);
  gmul2(166) <= to_unsigned(16#55#, 8);
  gmul2(167) <= to_unsigned(16#4B#, 8);
  gmul2(168) <= to_unsigned(16#49#, 8);
  gmul2(169) <= to_unsigned(16#4F#, 8);
  gmul2(170) <= to_unsigned(16#4D#, 8);
  gmul2(171) <= to_unsigned(16#43#, 8);
  gmul2(172) <= to_unsigned(16#41#, 8);
  gmul2(173) <= to_unsigned(16#47#, 8);
  gmul2(174) <= to_unsigned(16#45#, 8);
  gmul2(175) <= to_unsigned(16#7B#, 8);
  gmul2(176) <= to_unsigned(16#79#, 8);
  gmul2(177) <= to_unsigned(16#7F#, 8);
  gmul2(178) <= to_unsigned(16#7D#, 8);
  gmul2(179) <= to_unsigned(16#73#, 8);
  gmul2(180) <= to_unsigned(16#71#, 8);
  gmul2(181) <= to_unsigned(16#77#, 8);
  gmul2(182) <= to_unsigned(16#75#, 8);
  gmul2(183) <= to_unsigned(16#6B#, 8);
  gmul2(184) <= to_unsigned(16#69#, 8);
  gmul2(185) <= to_unsigned(16#6F#, 8);
  gmul2(186) <= to_unsigned(16#6D#, 8);
  gmul2(187) <= to_unsigned(16#63#, 8);
  gmul2(188) <= to_unsigned(16#61#, 8);
  gmul2(189) <= to_unsigned(16#67#, 8);
  gmul2(190) <= to_unsigned(16#65#, 8);
  gmul2(191) <= to_unsigned(16#9B#, 8);
  gmul2(192) <= to_unsigned(16#99#, 8);
  gmul2(193) <= to_unsigned(16#9F#, 8);
  gmul2(194) <= to_unsigned(16#9D#, 8);
  gmul2(195) <= to_unsigned(16#93#, 8);
  gmul2(196) <= to_unsigned(16#91#, 8);
  gmul2(197) <= to_unsigned(16#97#, 8);
  gmul2(198) <= to_unsigned(16#95#, 8);
  gmul2(199) <= to_unsigned(16#8B#, 8);
  gmul2(200) <= to_unsigned(16#89#, 8);
  gmul2(201) <= to_unsigned(16#8F#, 8);
  gmul2(202) <= to_unsigned(16#8D#, 8);
  gmul2(203) <= to_unsigned(16#83#, 8);
  gmul2(204) <= to_unsigned(16#81#, 8);
  gmul2(205) <= to_unsigned(16#87#, 8);
  gmul2(206) <= to_unsigned(16#85#, 8);
  gmul2(207) <= to_unsigned(16#BB#, 8);
  gmul2(208) <= to_unsigned(16#B9#, 8);
  gmul2(209) <= to_unsigned(16#BF#, 8);
  gmul2(210) <= to_unsigned(16#BD#, 8);
  gmul2(211) <= to_unsigned(16#B3#, 8);
  gmul2(212) <= to_unsigned(16#B1#, 8);
  gmul2(213) <= to_unsigned(16#B7#, 8);
  gmul2(214) <= to_unsigned(16#B5#, 8);
  gmul2(215) <= to_unsigned(16#AB#, 8);
  gmul2(216) <= to_unsigned(16#A9#, 8);
  gmul2(217) <= to_unsigned(16#AF#, 8);
  gmul2(218) <= to_unsigned(16#AD#, 8);
  gmul2(219) <= to_unsigned(16#A3#, 8);
  gmul2(220) <= to_unsigned(16#A1#, 8);
  gmul2(221) <= to_unsigned(16#A7#, 8);
  gmul2(222) <= to_unsigned(16#A5#, 8);
  gmul2(223) <= to_unsigned(16#DB#, 8);
  gmul2(224) <= to_unsigned(16#D9#, 8);
  gmul2(225) <= to_unsigned(16#DF#, 8);
  gmul2(226) <= to_unsigned(16#DD#, 8);
  gmul2(227) <= to_unsigned(16#D3#, 8);
  gmul2(228) <= to_unsigned(16#D1#, 8);
  gmul2(229) <= to_unsigned(16#D7#, 8);
  gmul2(230) <= to_unsigned(16#D5#, 8);
  gmul2(231) <= to_unsigned(16#CB#, 8);
  gmul2(232) <= to_unsigned(16#C9#, 8);
  gmul2(233) <= to_unsigned(16#CF#, 8);
  gmul2(234) <= to_unsigned(16#CD#, 8);
  gmul2(235) <= to_unsigned(16#C3#, 8);
  gmul2(236) <= to_unsigned(16#C1#, 8);
  gmul2(237) <= to_unsigned(16#C7#, 8);
  gmul2(238) <= to_unsigned(16#C5#, 8);
  gmul2(239) <= to_unsigned(16#FB#, 8);
  gmul2(240) <= to_unsigned(16#F9#, 8);
  gmul2(241) <= to_unsigned(16#FF#, 8);
  gmul2(242) <= to_unsigned(16#FD#, 8);
  gmul2(243) <= to_unsigned(16#F3#, 8);
  gmul2(244) <= to_unsigned(16#F1#, 8);
  gmul2(245) <= to_unsigned(16#F7#, 8);
  gmul2(246) <= to_unsigned(16#F5#, 8);
  gmul2(247) <= to_unsigned(16#EB#, 8);
  gmul2(248) <= to_unsigned(16#E9#, 8);
  gmul2(249) <= to_unsigned(16#EF#, 8);
  gmul2(250) <= to_unsigned(16#ED#, 8);
  gmul2(251) <= to_unsigned(16#E3#, 8);
  gmul2(252) <= to_unsigned(16#E1#, 8);
  gmul2(253) <= to_unsigned(16#E7#, 8);
  gmul2(254) <= to_unsigned(16#E5#, 8);
  gmul2(255) <= to_unsigned(16#E5#, 8);

  gmul3(0) <= to_unsigned(16#03#, 8);
  gmul3(1) <= to_unsigned(16#06#, 8);
  gmul3(2) <= to_unsigned(16#05#, 8);
  gmul3(3) <= to_unsigned(16#0C#, 8);
  gmul3(4) <= to_unsigned(16#0F#, 8);
  gmul3(5) <= to_unsigned(16#0A#, 8);
  gmul3(6) <= to_unsigned(16#09#, 8);
  gmul3(7) <= to_unsigned(16#18#, 8);
  gmul3(8) <= to_unsigned(16#1B#, 8);
  gmul3(9) <= to_unsigned(16#1E#, 8);
  gmul3(10) <= to_unsigned(16#1D#, 8);
  gmul3(11) <= to_unsigned(16#14#, 8);
  gmul3(12) <= to_unsigned(16#17#, 8);
  gmul3(13) <= to_unsigned(16#12#, 8);
  gmul3(14) <= to_unsigned(16#11#, 8);
  gmul3(15) <= to_unsigned(16#30#, 8);
  gmul3(16) <= to_unsigned(16#33#, 8);
  gmul3(17) <= to_unsigned(16#36#, 8);
  gmul3(18) <= to_unsigned(16#35#, 8);
  gmul3(19) <= to_unsigned(16#3C#, 8);
  gmul3(20) <= to_unsigned(16#3F#, 8);
  gmul3(21) <= to_unsigned(16#3A#, 8);
  gmul3(22) <= to_unsigned(16#39#, 8);
  gmul3(23) <= to_unsigned(16#28#, 8);
  gmul3(24) <= to_unsigned(16#2B#, 8);
  gmul3(25) <= to_unsigned(16#2E#, 8);
  gmul3(26) <= to_unsigned(16#2D#, 8);
  gmul3(27) <= to_unsigned(16#24#, 8);
  gmul3(28) <= to_unsigned(16#27#, 8);
  gmul3(29) <= to_unsigned(16#22#, 8);
  gmul3(30) <= to_unsigned(16#21#, 8);
  gmul3(31) <= to_unsigned(16#60#, 8);
  gmul3(32) <= to_unsigned(16#63#, 8);
  gmul3(33) <= to_unsigned(16#66#, 8);
  gmul3(34) <= to_unsigned(16#65#, 8);
  gmul3(35) <= to_unsigned(16#6C#, 8);
  gmul3(36) <= to_unsigned(16#6F#, 8);
  gmul3(37) <= to_unsigned(16#6A#, 8);
  gmul3(38) <= to_unsigned(16#69#, 8);
  gmul3(39) <= to_unsigned(16#78#, 8);
  gmul3(40) <= to_unsigned(16#7B#, 8);
  gmul3(41) <= to_unsigned(16#7E#, 8);
  gmul3(42) <= to_unsigned(16#7D#, 8);
  gmul3(43) <= to_unsigned(16#74#, 8);
  gmul3(44) <= to_unsigned(16#77#, 8);
  gmul3(45) <= to_unsigned(16#72#, 8);
  gmul3(46) <= to_unsigned(16#71#, 8);
  gmul3(47) <= to_unsigned(16#50#, 8);
  gmul3(48) <= to_unsigned(16#53#, 8);
  gmul3(49) <= to_unsigned(16#56#, 8);
  gmul3(50) <= to_unsigned(16#55#, 8);
  gmul3(51) <= to_unsigned(16#5C#, 8);
  gmul3(52) <= to_unsigned(16#5F#, 8);
  gmul3(53) <= to_unsigned(16#5A#, 8);
  gmul3(54) <= to_unsigned(16#59#, 8);
  gmul3(55) <= to_unsigned(16#48#, 8);
  gmul3(56) <= to_unsigned(16#4B#, 8);
  gmul3(57) <= to_unsigned(16#4E#, 8);
  gmul3(58) <= to_unsigned(16#4D#, 8);
  gmul3(59) <= to_unsigned(16#44#, 8);
  gmul3(60) <= to_unsigned(16#47#, 8);
  gmul3(61) <= to_unsigned(16#42#, 8);
  gmul3(62) <= to_unsigned(16#41#, 8);
  gmul3(63) <= to_unsigned(16#C0#, 8);
  gmul3(64) <= to_unsigned(16#C3#, 8);
  gmul3(65) <= to_unsigned(16#C6#, 8);
  gmul3(66) <= to_unsigned(16#C5#, 8);
  gmul3(67) <= to_unsigned(16#CC#, 8);
  gmul3(68) <= to_unsigned(16#CF#, 8);
  gmul3(69) <= to_unsigned(16#CA#, 8);
  gmul3(70) <= to_unsigned(16#C9#, 8);
  gmul3(71) <= to_unsigned(16#D8#, 8);
  gmul3(72) <= to_unsigned(16#DB#, 8);
  gmul3(73) <= to_unsigned(16#DE#, 8);
  gmul3(74) <= to_unsigned(16#DD#, 8);
  gmul3(75) <= to_unsigned(16#D4#, 8);
  gmul3(76) <= to_unsigned(16#D7#, 8);
  gmul3(77) <= to_unsigned(16#D2#, 8);
  gmul3(78) <= to_unsigned(16#D1#, 8);
  gmul3(79) <= to_unsigned(16#F0#, 8);
  gmul3(80) <= to_unsigned(16#F3#, 8);
  gmul3(81) <= to_unsigned(16#F6#, 8);
  gmul3(82) <= to_unsigned(16#F5#, 8);
  gmul3(83) <= to_unsigned(16#FC#, 8);
  gmul3(84) <= to_unsigned(16#FF#, 8);
  gmul3(85) <= to_unsigned(16#FA#, 8);
  gmul3(86) <= to_unsigned(16#F9#, 8);
  gmul3(87) <= to_unsigned(16#E8#, 8);
  gmul3(88) <= to_unsigned(16#EB#, 8);
  gmul3(89) <= to_unsigned(16#EE#, 8);
  gmul3(90) <= to_unsigned(16#ED#, 8);
  gmul3(91) <= to_unsigned(16#E4#, 8);
  gmul3(92) <= to_unsigned(16#E7#, 8);
  gmul3(93) <= to_unsigned(16#E2#, 8);
  gmul3(94) <= to_unsigned(16#E1#, 8);
  gmul3(95) <= to_unsigned(16#A0#, 8);
  gmul3(96) <= to_unsigned(16#A3#, 8);
  gmul3(97) <= to_unsigned(16#A6#, 8);
  gmul3(98) <= to_unsigned(16#A5#, 8);
  gmul3(99) <= to_unsigned(16#AC#, 8);
  gmul3(100) <= to_unsigned(16#AF#, 8);
  gmul3(101) <= to_unsigned(16#AA#, 8);
  gmul3(102) <= to_unsigned(16#A9#, 8);
  gmul3(103) <= to_unsigned(16#B8#, 8);
  gmul3(104) <= to_unsigned(16#BB#, 8);
  gmul3(105) <= to_unsigned(16#BE#, 8);
  gmul3(106) <= to_unsigned(16#BD#, 8);
  gmul3(107) <= to_unsigned(16#B4#, 8);
  gmul3(108) <= to_unsigned(16#B7#, 8);
  gmul3(109) <= to_unsigned(16#B2#, 8);
  gmul3(110) <= to_unsigned(16#B1#, 8);
  gmul3(111) <= to_unsigned(16#90#, 8);
  gmul3(112) <= to_unsigned(16#93#, 8);
  gmul3(113) <= to_unsigned(16#96#, 8);
  gmul3(114) <= to_unsigned(16#95#, 8);
  gmul3(115) <= to_unsigned(16#9C#, 8);
  gmul3(116) <= to_unsigned(16#9F#, 8);
  gmul3(117) <= to_unsigned(16#9A#, 8);
  gmul3(118) <= to_unsigned(16#99#, 8);
  gmul3(119) <= to_unsigned(16#88#, 8);
  gmul3(120) <= to_unsigned(16#8B#, 8);
  gmul3(121) <= to_unsigned(16#8E#, 8);
  gmul3(122) <= to_unsigned(16#8D#, 8);
  gmul3(123) <= to_unsigned(16#84#, 8);
  gmul3(124) <= to_unsigned(16#87#, 8);
  gmul3(125) <= to_unsigned(16#82#, 8);
  gmul3(126) <= to_unsigned(16#81#, 8);
  gmul3(127) <= to_unsigned(16#9B#, 8);
  gmul3(128) <= to_unsigned(16#98#, 8);
  gmul3(129) <= to_unsigned(16#9D#, 8);
  gmul3(130) <= to_unsigned(16#9E#, 8);
  gmul3(131) <= to_unsigned(16#97#, 8);
  gmul3(132) <= to_unsigned(16#94#, 8);
  gmul3(133) <= to_unsigned(16#91#, 8);
  gmul3(134) <= to_unsigned(16#92#, 8);
  gmul3(135) <= to_unsigned(16#83#, 8);
  gmul3(136) <= to_unsigned(16#80#, 8);
  gmul3(137) <= to_unsigned(16#85#, 8);
  gmul3(138) <= to_unsigned(16#86#, 8);
  gmul3(139) <= to_unsigned(16#8F#, 8);
  gmul3(140) <= to_unsigned(16#8C#, 8);
  gmul3(141) <= to_unsigned(16#89#, 8);
  gmul3(142) <= to_unsigned(16#8A#, 8);
  gmul3(143) <= to_unsigned(16#AB#, 8);
  gmul3(144) <= to_unsigned(16#A8#, 8);
  gmul3(145) <= to_unsigned(16#AD#, 8);
  gmul3(146) <= to_unsigned(16#AE#, 8);
  gmul3(147) <= to_unsigned(16#A7#, 8);
  gmul3(148) <= to_unsigned(16#A4#, 8);
  gmul3(149) <= to_unsigned(16#A1#, 8);
  gmul3(150) <= to_unsigned(16#A2#, 8);
  gmul3(151) <= to_unsigned(16#B3#, 8);
  gmul3(152) <= to_unsigned(16#B0#, 8);
  gmul3(153) <= to_unsigned(16#B5#, 8);
  gmul3(154) <= to_unsigned(16#B6#, 8);
  gmul3(155) <= to_unsigned(16#BF#, 8);
  gmul3(156) <= to_unsigned(16#BC#, 8);
  gmul3(157) <= to_unsigned(16#B9#, 8);
  gmul3(158) <= to_unsigned(16#BA#, 8);
  gmul3(159) <= to_unsigned(16#FB#, 8);
  gmul3(160) <= to_unsigned(16#F8#, 8);
  gmul3(161) <= to_unsigned(16#FD#, 8);
  gmul3(162) <= to_unsigned(16#FE#, 8);
  gmul3(163) <= to_unsigned(16#F7#, 8);
  gmul3(164) <= to_unsigned(16#F4#, 8);
  gmul3(165) <= to_unsigned(16#F1#, 8);
  gmul3(166) <= to_unsigned(16#F2#, 8);
  gmul3(167) <= to_unsigned(16#E3#, 8);
  gmul3(168) <= to_unsigned(16#E0#, 8);
  gmul3(169) <= to_unsigned(16#E5#, 8);
  gmul3(170) <= to_unsigned(16#E6#, 8);
  gmul3(171) <= to_unsigned(16#EF#, 8);
  gmul3(172) <= to_unsigned(16#EC#, 8);
  gmul3(173) <= to_unsigned(16#E9#, 8);
  gmul3(174) <= to_unsigned(16#EA#, 8);
  gmul3(175) <= to_unsigned(16#CB#, 8);
  gmul3(176) <= to_unsigned(16#C8#, 8);
  gmul3(177) <= to_unsigned(16#CD#, 8);
  gmul3(178) <= to_unsigned(16#CE#, 8);
  gmul3(179) <= to_unsigned(16#C7#, 8);
  gmul3(180) <= to_unsigned(16#C4#, 8);
  gmul3(181) <= to_unsigned(16#C1#, 8);
  gmul3(182) <= to_unsigned(16#C2#, 8);
  gmul3(183) <= to_unsigned(16#D3#, 8);
  gmul3(184) <= to_unsigned(16#D0#, 8);
  gmul3(185) <= to_unsigned(16#D5#, 8);
  gmul3(186) <= to_unsigned(16#D6#, 8);
  gmul3(187) <= to_unsigned(16#DF#, 8);
  gmul3(188) <= to_unsigned(16#DC#, 8);
  gmul3(189) <= to_unsigned(16#D9#, 8);
  gmul3(190) <= to_unsigned(16#DA#, 8);
  gmul3(191) <= to_unsigned(16#5B#, 8);
  gmul3(192) <= to_unsigned(16#58#, 8);
  gmul3(193) <= to_unsigned(16#5D#, 8);
  gmul3(194) <= to_unsigned(16#5E#, 8);
  gmul3(195) <= to_unsigned(16#57#, 8);
  gmul3(196) <= to_unsigned(16#54#, 8);
  gmul3(197) <= to_unsigned(16#51#, 8);
  gmul3(198) <= to_unsigned(16#52#, 8);
  gmul3(199) <= to_unsigned(16#43#, 8);
  gmul3(200) <= to_unsigned(16#40#, 8);
  gmul3(201) <= to_unsigned(16#45#, 8);
  gmul3(202) <= to_unsigned(16#46#, 8);
  gmul3(203) <= to_unsigned(16#4F#, 8);
  gmul3(204) <= to_unsigned(16#4C#, 8);
  gmul3(205) <= to_unsigned(16#49#, 8);
  gmul3(206) <= to_unsigned(16#4A#, 8);
  gmul3(207) <= to_unsigned(16#6B#, 8);
  gmul3(208) <= to_unsigned(16#68#, 8);
  gmul3(209) <= to_unsigned(16#6D#, 8);
  gmul3(210) <= to_unsigned(16#6E#, 8);
  gmul3(211) <= to_unsigned(16#67#, 8);
  gmul3(212) <= to_unsigned(16#64#, 8);
  gmul3(213) <= to_unsigned(16#61#, 8);
  gmul3(214) <= to_unsigned(16#62#, 8);
  gmul3(215) <= to_unsigned(16#73#, 8);
  gmul3(216) <= to_unsigned(16#70#, 8);
  gmul3(217) <= to_unsigned(16#75#, 8);
  gmul3(218) <= to_unsigned(16#76#, 8);
  gmul3(219) <= to_unsigned(16#7F#, 8);
  gmul3(220) <= to_unsigned(16#7C#, 8);
  gmul3(221) <= to_unsigned(16#79#, 8);
  gmul3(222) <= to_unsigned(16#7A#, 8);
  gmul3(223) <= to_unsigned(16#3B#, 8);
  gmul3(224) <= to_unsigned(16#38#, 8);
  gmul3(225) <= to_unsigned(16#3D#, 8);
  gmul3(226) <= to_unsigned(16#3E#, 8);
  gmul3(227) <= to_unsigned(16#37#, 8);
  gmul3(228) <= to_unsigned(16#34#, 8);
  gmul3(229) <= to_unsigned(16#31#, 8);
  gmul3(230) <= to_unsigned(16#32#, 8);
  gmul3(231) <= to_unsigned(16#23#, 8);
  gmul3(232) <= to_unsigned(16#20#, 8);
  gmul3(233) <= to_unsigned(16#25#, 8);
  gmul3(234) <= to_unsigned(16#26#, 8);
  gmul3(235) <= to_unsigned(16#2F#, 8);
  gmul3(236) <= to_unsigned(16#2C#, 8);
  gmul3(237) <= to_unsigned(16#29#, 8);
  gmul3(238) <= to_unsigned(16#2A#, 8);
  gmul3(239) <= to_unsigned(16#0B#, 8);
  gmul3(240) <= to_unsigned(16#08#, 8);
  gmul3(241) <= to_unsigned(16#0D#, 8);
  gmul3(242) <= to_unsigned(16#0E#, 8);
  gmul3(243) <= to_unsigned(16#07#, 8);
  gmul3(244) <= to_unsigned(16#04#, 8);
  gmul3(245) <= to_unsigned(16#01#, 8);
  gmul3(246) <= to_unsigned(16#02#, 8);
  gmul3(247) <= to_unsigned(16#13#, 8);
  gmul3(248) <= to_unsigned(16#10#, 8);
  gmul3(249) <= to_unsigned(16#15#, 8);
  gmul3(250) <= to_unsigned(16#16#, 8);
  gmul3(251) <= to_unsigned(16#1F#, 8);
  gmul3(252) <= to_unsigned(16#1C#, 8);
  gmul3(253) <= to_unsigned(16#19#, 8);
  gmul3(254) <= to_unsigned(16#1A#, 8);
  gmul3(255) <= to_unsigned(16#1A#, 8);

  gmul2_1(0) <= to_unsigned(16#02#, 8);
  gmul2_1(1) <= to_unsigned(16#04#, 8);
  gmul2_1(2) <= to_unsigned(16#06#, 8);
  gmul2_1(3) <= to_unsigned(16#08#, 8);
  gmul2_1(4) <= to_unsigned(16#0A#, 8);
  gmul2_1(5) <= to_unsigned(16#0C#, 8);
  gmul2_1(6) <= to_unsigned(16#0E#, 8);
  gmul2_1(7) <= to_unsigned(16#10#, 8);
  gmul2_1(8) <= to_unsigned(16#12#, 8);
  gmul2_1(9) <= to_unsigned(16#14#, 8);
  gmul2_1(10) <= to_unsigned(16#16#, 8);
  gmul2_1(11) <= to_unsigned(16#18#, 8);
  gmul2_1(12) <= to_unsigned(16#1A#, 8);
  gmul2_1(13) <= to_unsigned(16#1C#, 8);
  gmul2_1(14) <= to_unsigned(16#1E#, 8);
  gmul2_1(15) <= to_unsigned(16#20#, 8);
  gmul2_1(16) <= to_unsigned(16#22#, 8);
  gmul2_1(17) <= to_unsigned(16#24#, 8);
  gmul2_1(18) <= to_unsigned(16#26#, 8);
  gmul2_1(19) <= to_unsigned(16#28#, 8);
  gmul2_1(20) <= to_unsigned(16#2A#, 8);
  gmul2_1(21) <= to_unsigned(16#2C#, 8);
  gmul2_1(22) <= to_unsigned(16#2E#, 8);
  gmul2_1(23) <= to_unsigned(16#30#, 8);
  gmul2_1(24) <= to_unsigned(16#32#, 8);
  gmul2_1(25) <= to_unsigned(16#34#, 8);
  gmul2_1(26) <= to_unsigned(16#36#, 8);
  gmul2_1(27) <= to_unsigned(16#38#, 8);
  gmul2_1(28) <= to_unsigned(16#3A#, 8);
  gmul2_1(29) <= to_unsigned(16#3C#, 8);
  gmul2_1(30) <= to_unsigned(16#3E#, 8);
  gmul2_1(31) <= to_unsigned(16#40#, 8);
  gmul2_1(32) <= to_unsigned(16#42#, 8);
  gmul2_1(33) <= to_unsigned(16#44#, 8);
  gmul2_1(34) <= to_unsigned(16#46#, 8);
  gmul2_1(35) <= to_unsigned(16#48#, 8);
  gmul2_1(36) <= to_unsigned(16#4A#, 8);
  gmul2_1(37) <= to_unsigned(16#4C#, 8);
  gmul2_1(38) <= to_unsigned(16#4E#, 8);
  gmul2_1(39) <= to_unsigned(16#50#, 8);
  gmul2_1(40) <= to_unsigned(16#52#, 8);
  gmul2_1(41) <= to_unsigned(16#54#, 8);
  gmul2_1(42) <= to_unsigned(16#56#, 8);
  gmul2_1(43) <= to_unsigned(16#58#, 8);
  gmul2_1(44) <= to_unsigned(16#5A#, 8);
  gmul2_1(45) <= to_unsigned(16#5C#, 8);
  gmul2_1(46) <= to_unsigned(16#5E#, 8);
  gmul2_1(47) <= to_unsigned(16#60#, 8);
  gmul2_1(48) <= to_unsigned(16#62#, 8);
  gmul2_1(49) <= to_unsigned(16#64#, 8);
  gmul2_1(50) <= to_unsigned(16#66#, 8);
  gmul2_1(51) <= to_unsigned(16#68#, 8);
  gmul2_1(52) <= to_unsigned(16#6A#, 8);
  gmul2_1(53) <= to_unsigned(16#6C#, 8);
  gmul2_1(54) <= to_unsigned(16#6E#, 8);
  gmul2_1(55) <= to_unsigned(16#70#, 8);
  gmul2_1(56) <= to_unsigned(16#72#, 8);
  gmul2_1(57) <= to_unsigned(16#74#, 8);
  gmul2_1(58) <= to_unsigned(16#76#, 8);
  gmul2_1(59) <= to_unsigned(16#78#, 8);
  gmul2_1(60) <= to_unsigned(16#7A#, 8);
  gmul2_1(61) <= to_unsigned(16#7C#, 8);
  gmul2_1(62) <= to_unsigned(16#7E#, 8);
  gmul2_1(63) <= to_unsigned(16#80#, 8);
  gmul2_1(64) <= to_unsigned(16#82#, 8);
  gmul2_1(65) <= to_unsigned(16#84#, 8);
  gmul2_1(66) <= to_unsigned(16#86#, 8);
  gmul2_1(67) <= to_unsigned(16#88#, 8);
  gmul2_1(68) <= to_unsigned(16#8A#, 8);
  gmul2_1(69) <= to_unsigned(16#8C#, 8);
  gmul2_1(70) <= to_unsigned(16#8E#, 8);
  gmul2_1(71) <= to_unsigned(16#90#, 8);
  gmul2_1(72) <= to_unsigned(16#92#, 8);
  gmul2_1(73) <= to_unsigned(16#94#, 8);
  gmul2_1(74) <= to_unsigned(16#96#, 8);
  gmul2_1(75) <= to_unsigned(16#98#, 8);
  gmul2_1(76) <= to_unsigned(16#9A#, 8);
  gmul2_1(77) <= to_unsigned(16#9C#, 8);
  gmul2_1(78) <= to_unsigned(16#9E#, 8);
  gmul2_1(79) <= to_unsigned(16#A0#, 8);
  gmul2_1(80) <= to_unsigned(16#A2#, 8);
  gmul2_1(81) <= to_unsigned(16#A4#, 8);
  gmul2_1(82) <= to_unsigned(16#A6#, 8);
  gmul2_1(83) <= to_unsigned(16#A8#, 8);
  gmul2_1(84) <= to_unsigned(16#AA#, 8);
  gmul2_1(85) <= to_unsigned(16#AC#, 8);
  gmul2_1(86) <= to_unsigned(16#AE#, 8);
  gmul2_1(87) <= to_unsigned(16#B0#, 8);
  gmul2_1(88) <= to_unsigned(16#B2#, 8);
  gmul2_1(89) <= to_unsigned(16#B4#, 8);
  gmul2_1(90) <= to_unsigned(16#B6#, 8);
  gmul2_1(91) <= to_unsigned(16#B8#, 8);
  gmul2_1(92) <= to_unsigned(16#BA#, 8);
  gmul2_1(93) <= to_unsigned(16#BC#, 8);
  gmul2_1(94) <= to_unsigned(16#BE#, 8);
  gmul2_1(95) <= to_unsigned(16#C0#, 8);
  gmul2_1(96) <= to_unsigned(16#C2#, 8);
  gmul2_1(97) <= to_unsigned(16#C4#, 8);
  gmul2_1(98) <= to_unsigned(16#C6#, 8);
  gmul2_1(99) <= to_unsigned(16#C8#, 8);
  gmul2_1(100) <= to_unsigned(16#CA#, 8);
  gmul2_1(101) <= to_unsigned(16#CC#, 8);
  gmul2_1(102) <= to_unsigned(16#CE#, 8);
  gmul2_1(103) <= to_unsigned(16#D0#, 8);
  gmul2_1(104) <= to_unsigned(16#D2#, 8);
  gmul2_1(105) <= to_unsigned(16#D4#, 8);
  gmul2_1(106) <= to_unsigned(16#D6#, 8);
  gmul2_1(107) <= to_unsigned(16#D8#, 8);
  gmul2_1(108) <= to_unsigned(16#DA#, 8);
  gmul2_1(109) <= to_unsigned(16#DC#, 8);
  gmul2_1(110) <= to_unsigned(16#DE#, 8);
  gmul2_1(111) <= to_unsigned(16#E0#, 8);
  gmul2_1(112) <= to_unsigned(16#E2#, 8);
  gmul2_1(113) <= to_unsigned(16#E4#, 8);
  gmul2_1(114) <= to_unsigned(16#E6#, 8);
  gmul2_1(115) <= to_unsigned(16#E8#, 8);
  gmul2_1(116) <= to_unsigned(16#EA#, 8);
  gmul2_1(117) <= to_unsigned(16#EC#, 8);
  gmul2_1(118) <= to_unsigned(16#EE#, 8);
  gmul2_1(119) <= to_unsigned(16#F0#, 8);
  gmul2_1(120) <= to_unsigned(16#F2#, 8);
  gmul2_1(121) <= to_unsigned(16#F4#, 8);
  gmul2_1(122) <= to_unsigned(16#F6#, 8);
  gmul2_1(123) <= to_unsigned(16#F8#, 8);
  gmul2_1(124) <= to_unsigned(16#FA#, 8);
  gmul2_1(125) <= to_unsigned(16#FC#, 8);
  gmul2_1(126) <= to_unsigned(16#FE#, 8);
  gmul2_1(127) <= to_unsigned(16#1B#, 8);
  gmul2_1(128) <= to_unsigned(16#19#, 8);
  gmul2_1(129) <= to_unsigned(16#1F#, 8);
  gmul2_1(130) <= to_unsigned(16#1D#, 8);
  gmul2_1(131) <= to_unsigned(16#13#, 8);
  gmul2_1(132) <= to_unsigned(16#11#, 8);
  gmul2_1(133) <= to_unsigned(16#17#, 8);
  gmul2_1(134) <= to_unsigned(16#15#, 8);
  gmul2_1(135) <= to_unsigned(16#0B#, 8);
  gmul2_1(136) <= to_unsigned(16#09#, 8);
  gmul2_1(137) <= to_unsigned(16#0F#, 8);
  gmul2_1(138) <= to_unsigned(16#0D#, 8);
  gmul2_1(139) <= to_unsigned(16#03#, 8);
  gmul2_1(140) <= to_unsigned(16#01#, 8);
  gmul2_1(141) <= to_unsigned(16#07#, 8);
  gmul2_1(142) <= to_unsigned(16#05#, 8);
  gmul2_1(143) <= to_unsigned(16#3B#, 8);
  gmul2_1(144) <= to_unsigned(16#39#, 8);
  gmul2_1(145) <= to_unsigned(16#3F#, 8);
  gmul2_1(146) <= to_unsigned(16#3D#, 8);
  gmul2_1(147) <= to_unsigned(16#33#, 8);
  gmul2_1(148) <= to_unsigned(16#31#, 8);
  gmul2_1(149) <= to_unsigned(16#37#, 8);
  gmul2_1(150) <= to_unsigned(16#35#, 8);
  gmul2_1(151) <= to_unsigned(16#2B#, 8);
  gmul2_1(152) <= to_unsigned(16#29#, 8);
  gmul2_1(153) <= to_unsigned(16#2F#, 8);
  gmul2_1(154) <= to_unsigned(16#2D#, 8);
  gmul2_1(155) <= to_unsigned(16#23#, 8);
  gmul2_1(156) <= to_unsigned(16#21#, 8);
  gmul2_1(157) <= to_unsigned(16#27#, 8);
  gmul2_1(158) <= to_unsigned(16#25#, 8);
  gmul2_1(159) <= to_unsigned(16#5B#, 8);
  gmul2_1(160) <= to_unsigned(16#59#, 8);
  gmul2_1(161) <= to_unsigned(16#5F#, 8);
  gmul2_1(162) <= to_unsigned(16#5D#, 8);
  gmul2_1(163) <= to_unsigned(16#53#, 8);
  gmul2_1(164) <= to_unsigned(16#51#, 8);
  gmul2_1(165) <= to_unsigned(16#57#, 8);
  gmul2_1(166) <= to_unsigned(16#55#, 8);
  gmul2_1(167) <= to_unsigned(16#4B#, 8);
  gmul2_1(168) <= to_unsigned(16#49#, 8);
  gmul2_1(169) <= to_unsigned(16#4F#, 8);
  gmul2_1(170) <= to_unsigned(16#4D#, 8);
  gmul2_1(171) <= to_unsigned(16#43#, 8);
  gmul2_1(172) <= to_unsigned(16#41#, 8);
  gmul2_1(173) <= to_unsigned(16#47#, 8);
  gmul2_1(174) <= to_unsigned(16#45#, 8);
  gmul2_1(175) <= to_unsigned(16#7B#, 8);
  gmul2_1(176) <= to_unsigned(16#79#, 8);
  gmul2_1(177) <= to_unsigned(16#7F#, 8);
  gmul2_1(178) <= to_unsigned(16#7D#, 8);
  gmul2_1(179) <= to_unsigned(16#73#, 8);
  gmul2_1(180) <= to_unsigned(16#71#, 8);
  gmul2_1(181) <= to_unsigned(16#77#, 8);
  gmul2_1(182) <= to_unsigned(16#75#, 8);
  gmul2_1(183) <= to_unsigned(16#6B#, 8);
  gmul2_1(184) <= to_unsigned(16#69#, 8);
  gmul2_1(185) <= to_unsigned(16#6F#, 8);
  gmul2_1(186) <= to_unsigned(16#6D#, 8);
  gmul2_1(187) <= to_unsigned(16#63#, 8);
  gmul2_1(188) <= to_unsigned(16#61#, 8);
  gmul2_1(189) <= to_unsigned(16#67#, 8);
  gmul2_1(190) <= to_unsigned(16#65#, 8);
  gmul2_1(191) <= to_unsigned(16#9B#, 8);
  gmul2_1(192) <= to_unsigned(16#99#, 8);
  gmul2_1(193) <= to_unsigned(16#9F#, 8);
  gmul2_1(194) <= to_unsigned(16#9D#, 8);
  gmul2_1(195) <= to_unsigned(16#93#, 8);
  gmul2_1(196) <= to_unsigned(16#91#, 8);
  gmul2_1(197) <= to_unsigned(16#97#, 8);
  gmul2_1(198) <= to_unsigned(16#95#, 8);
  gmul2_1(199) <= to_unsigned(16#8B#, 8);
  gmul2_1(200) <= to_unsigned(16#89#, 8);
  gmul2_1(201) <= to_unsigned(16#8F#, 8);
  gmul2_1(202) <= to_unsigned(16#8D#, 8);
  gmul2_1(203) <= to_unsigned(16#83#, 8);
  gmul2_1(204) <= to_unsigned(16#81#, 8);
  gmul2_1(205) <= to_unsigned(16#87#, 8);
  gmul2_1(206) <= to_unsigned(16#85#, 8);
  gmul2_1(207) <= to_unsigned(16#BB#, 8);
  gmul2_1(208) <= to_unsigned(16#B9#, 8);
  gmul2_1(209) <= to_unsigned(16#BF#, 8);
  gmul2_1(210) <= to_unsigned(16#BD#, 8);
  gmul2_1(211) <= to_unsigned(16#B3#, 8);
  gmul2_1(212) <= to_unsigned(16#B1#, 8);
  gmul2_1(213) <= to_unsigned(16#B7#, 8);
  gmul2_1(214) <= to_unsigned(16#B5#, 8);
  gmul2_1(215) <= to_unsigned(16#AB#, 8);
  gmul2_1(216) <= to_unsigned(16#A9#, 8);
  gmul2_1(217) <= to_unsigned(16#AF#, 8);
  gmul2_1(218) <= to_unsigned(16#AD#, 8);
  gmul2_1(219) <= to_unsigned(16#A3#, 8);
  gmul2_1(220) <= to_unsigned(16#A1#, 8);
  gmul2_1(221) <= to_unsigned(16#A7#, 8);
  gmul2_1(222) <= to_unsigned(16#A5#, 8);
  gmul2_1(223) <= to_unsigned(16#DB#, 8);
  gmul2_1(224) <= to_unsigned(16#D9#, 8);
  gmul2_1(225) <= to_unsigned(16#DF#, 8);
  gmul2_1(226) <= to_unsigned(16#DD#, 8);
  gmul2_1(227) <= to_unsigned(16#D3#, 8);
  gmul2_1(228) <= to_unsigned(16#D1#, 8);
  gmul2_1(229) <= to_unsigned(16#D7#, 8);
  gmul2_1(230) <= to_unsigned(16#D5#, 8);
  gmul2_1(231) <= to_unsigned(16#CB#, 8);
  gmul2_1(232) <= to_unsigned(16#C9#, 8);
  gmul2_1(233) <= to_unsigned(16#CF#, 8);
  gmul2_1(234) <= to_unsigned(16#CD#, 8);
  gmul2_1(235) <= to_unsigned(16#C3#, 8);
  gmul2_1(236) <= to_unsigned(16#C1#, 8);
  gmul2_1(237) <= to_unsigned(16#C7#, 8);
  gmul2_1(238) <= to_unsigned(16#C5#, 8);
  gmul2_1(239) <= to_unsigned(16#FB#, 8);
  gmul2_1(240) <= to_unsigned(16#F9#, 8);
  gmul2_1(241) <= to_unsigned(16#FF#, 8);
  gmul2_1(242) <= to_unsigned(16#FD#, 8);
  gmul2_1(243) <= to_unsigned(16#F3#, 8);
  gmul2_1(244) <= to_unsigned(16#F1#, 8);
  gmul2_1(245) <= to_unsigned(16#F7#, 8);
  gmul2_1(246) <= to_unsigned(16#F5#, 8);
  gmul2_1(247) <= to_unsigned(16#EB#, 8);
  gmul2_1(248) <= to_unsigned(16#E9#, 8);
  gmul2_1(249) <= to_unsigned(16#EF#, 8);
  gmul2_1(250) <= to_unsigned(16#ED#, 8);
  gmul2_1(251) <= to_unsigned(16#E3#, 8);
  gmul2_1(252) <= to_unsigned(16#E1#, 8);
  gmul2_1(253) <= to_unsigned(16#E7#, 8);
  gmul2_1(254) <= to_unsigned(16#E5#, 8);
  gmul2_1(255) <= to_unsigned(16#E5#, 8);

  gmul3_1(0) <= to_unsigned(16#03#, 8);
  gmul3_1(1) <= to_unsigned(16#06#, 8);
  gmul3_1(2) <= to_unsigned(16#05#, 8);
  gmul3_1(3) <= to_unsigned(16#0C#, 8);
  gmul3_1(4) <= to_unsigned(16#0F#, 8);
  gmul3_1(5) <= to_unsigned(16#0A#, 8);
  gmul3_1(6) <= to_unsigned(16#09#, 8);
  gmul3_1(7) <= to_unsigned(16#18#, 8);
  gmul3_1(8) <= to_unsigned(16#1B#, 8);
  gmul3_1(9) <= to_unsigned(16#1E#, 8);
  gmul3_1(10) <= to_unsigned(16#1D#, 8);
  gmul3_1(11) <= to_unsigned(16#14#, 8);
  gmul3_1(12) <= to_unsigned(16#17#, 8);
  gmul3_1(13) <= to_unsigned(16#12#, 8);
  gmul3_1(14) <= to_unsigned(16#11#, 8);
  gmul3_1(15) <= to_unsigned(16#30#, 8);
  gmul3_1(16) <= to_unsigned(16#33#, 8);
  gmul3_1(17) <= to_unsigned(16#36#, 8);
  gmul3_1(18) <= to_unsigned(16#35#, 8);
  gmul3_1(19) <= to_unsigned(16#3C#, 8);
  gmul3_1(20) <= to_unsigned(16#3F#, 8);
  gmul3_1(21) <= to_unsigned(16#3A#, 8);
  gmul3_1(22) <= to_unsigned(16#39#, 8);
  gmul3_1(23) <= to_unsigned(16#28#, 8);
  gmul3_1(24) <= to_unsigned(16#2B#, 8);
  gmul3_1(25) <= to_unsigned(16#2E#, 8);
  gmul3_1(26) <= to_unsigned(16#2D#, 8);
  gmul3_1(27) <= to_unsigned(16#24#, 8);
  gmul3_1(28) <= to_unsigned(16#27#, 8);
  gmul3_1(29) <= to_unsigned(16#22#, 8);
  gmul3_1(30) <= to_unsigned(16#21#, 8);
  gmul3_1(31) <= to_unsigned(16#60#, 8);
  gmul3_1(32) <= to_unsigned(16#63#, 8);
  gmul3_1(33) <= to_unsigned(16#66#, 8);
  gmul3_1(34) <= to_unsigned(16#65#, 8);
  gmul3_1(35) <= to_unsigned(16#6C#, 8);
  gmul3_1(36) <= to_unsigned(16#6F#, 8);
  gmul3_1(37) <= to_unsigned(16#6A#, 8);
  gmul3_1(38) <= to_unsigned(16#69#, 8);
  gmul3_1(39) <= to_unsigned(16#78#, 8);
  gmul3_1(40) <= to_unsigned(16#7B#, 8);
  gmul3_1(41) <= to_unsigned(16#7E#, 8);
  gmul3_1(42) <= to_unsigned(16#7D#, 8);
  gmul3_1(43) <= to_unsigned(16#74#, 8);
  gmul3_1(44) <= to_unsigned(16#77#, 8);
  gmul3_1(45) <= to_unsigned(16#72#, 8);
  gmul3_1(46) <= to_unsigned(16#71#, 8);
  gmul3_1(47) <= to_unsigned(16#50#, 8);
  gmul3_1(48) <= to_unsigned(16#53#, 8);
  gmul3_1(49) <= to_unsigned(16#56#, 8);
  gmul3_1(50) <= to_unsigned(16#55#, 8);
  gmul3_1(51) <= to_unsigned(16#5C#, 8);
  gmul3_1(52) <= to_unsigned(16#5F#, 8);
  gmul3_1(53) <= to_unsigned(16#5A#, 8);
  gmul3_1(54) <= to_unsigned(16#59#, 8);
  gmul3_1(55) <= to_unsigned(16#48#, 8);
  gmul3_1(56) <= to_unsigned(16#4B#, 8);
  gmul3_1(57) <= to_unsigned(16#4E#, 8);
  gmul3_1(58) <= to_unsigned(16#4D#, 8);
  gmul3_1(59) <= to_unsigned(16#44#, 8);
  gmul3_1(60) <= to_unsigned(16#47#, 8);
  gmul3_1(61) <= to_unsigned(16#42#, 8);
  gmul3_1(62) <= to_unsigned(16#41#, 8);
  gmul3_1(63) <= to_unsigned(16#C0#, 8);
  gmul3_1(64) <= to_unsigned(16#C3#, 8);
  gmul3_1(65) <= to_unsigned(16#C6#, 8);
  gmul3_1(66) <= to_unsigned(16#C5#, 8);
  gmul3_1(67) <= to_unsigned(16#CC#, 8);
  gmul3_1(68) <= to_unsigned(16#CF#, 8);
  gmul3_1(69) <= to_unsigned(16#CA#, 8);
  gmul3_1(70) <= to_unsigned(16#C9#, 8);
  gmul3_1(71) <= to_unsigned(16#D8#, 8);
  gmul3_1(72) <= to_unsigned(16#DB#, 8);
  gmul3_1(73) <= to_unsigned(16#DE#, 8);
  gmul3_1(74) <= to_unsigned(16#DD#, 8);
  gmul3_1(75) <= to_unsigned(16#D4#, 8);
  gmul3_1(76) <= to_unsigned(16#D7#, 8);
  gmul3_1(77) <= to_unsigned(16#D2#, 8);
  gmul3_1(78) <= to_unsigned(16#D1#, 8);
  gmul3_1(79) <= to_unsigned(16#F0#, 8);
  gmul3_1(80) <= to_unsigned(16#F3#, 8);
  gmul3_1(81) <= to_unsigned(16#F6#, 8);
  gmul3_1(82) <= to_unsigned(16#F5#, 8);
  gmul3_1(83) <= to_unsigned(16#FC#, 8);
  gmul3_1(84) <= to_unsigned(16#FF#, 8);
  gmul3_1(85) <= to_unsigned(16#FA#, 8);
  gmul3_1(86) <= to_unsigned(16#F9#, 8);
  gmul3_1(87) <= to_unsigned(16#E8#, 8);
  gmul3_1(88) <= to_unsigned(16#EB#, 8);
  gmul3_1(89) <= to_unsigned(16#EE#, 8);
  gmul3_1(90) <= to_unsigned(16#ED#, 8);
  gmul3_1(91) <= to_unsigned(16#E4#, 8);
  gmul3_1(92) <= to_unsigned(16#E7#, 8);
  gmul3_1(93) <= to_unsigned(16#E2#, 8);
  gmul3_1(94) <= to_unsigned(16#E1#, 8);
  gmul3_1(95) <= to_unsigned(16#A0#, 8);
  gmul3_1(96) <= to_unsigned(16#A3#, 8);
  gmul3_1(97) <= to_unsigned(16#A6#, 8);
  gmul3_1(98) <= to_unsigned(16#A5#, 8);
  gmul3_1(99) <= to_unsigned(16#AC#, 8);
  gmul3_1(100) <= to_unsigned(16#AF#, 8);
  gmul3_1(101) <= to_unsigned(16#AA#, 8);
  gmul3_1(102) <= to_unsigned(16#A9#, 8);
  gmul3_1(103) <= to_unsigned(16#B8#, 8);
  gmul3_1(104) <= to_unsigned(16#BB#, 8);
  gmul3_1(105) <= to_unsigned(16#BE#, 8);
  gmul3_1(106) <= to_unsigned(16#BD#, 8);
  gmul3_1(107) <= to_unsigned(16#B4#, 8);
  gmul3_1(108) <= to_unsigned(16#B7#, 8);
  gmul3_1(109) <= to_unsigned(16#B2#, 8);
  gmul3_1(110) <= to_unsigned(16#B1#, 8);
  gmul3_1(111) <= to_unsigned(16#90#, 8);
  gmul3_1(112) <= to_unsigned(16#93#, 8);
  gmul3_1(113) <= to_unsigned(16#96#, 8);
  gmul3_1(114) <= to_unsigned(16#95#, 8);
  gmul3_1(115) <= to_unsigned(16#9C#, 8);
  gmul3_1(116) <= to_unsigned(16#9F#, 8);
  gmul3_1(117) <= to_unsigned(16#9A#, 8);
  gmul3_1(118) <= to_unsigned(16#99#, 8);
  gmul3_1(119) <= to_unsigned(16#88#, 8);
  gmul3_1(120) <= to_unsigned(16#8B#, 8);
  gmul3_1(121) <= to_unsigned(16#8E#, 8);
  gmul3_1(122) <= to_unsigned(16#8D#, 8);
  gmul3_1(123) <= to_unsigned(16#84#, 8);
  gmul3_1(124) <= to_unsigned(16#87#, 8);
  gmul3_1(125) <= to_unsigned(16#82#, 8);
  gmul3_1(126) <= to_unsigned(16#81#, 8);
  gmul3_1(127) <= to_unsigned(16#9B#, 8);
  gmul3_1(128) <= to_unsigned(16#98#, 8);
  gmul3_1(129) <= to_unsigned(16#9D#, 8);
  gmul3_1(130) <= to_unsigned(16#9E#, 8);
  gmul3_1(131) <= to_unsigned(16#97#, 8);
  gmul3_1(132) <= to_unsigned(16#94#, 8);
  gmul3_1(133) <= to_unsigned(16#91#, 8);
  gmul3_1(134) <= to_unsigned(16#92#, 8);
  gmul3_1(135) <= to_unsigned(16#83#, 8);
  gmul3_1(136) <= to_unsigned(16#80#, 8);
  gmul3_1(137) <= to_unsigned(16#85#, 8);
  gmul3_1(138) <= to_unsigned(16#86#, 8);
  gmul3_1(139) <= to_unsigned(16#8F#, 8);
  gmul3_1(140) <= to_unsigned(16#8C#, 8);
  gmul3_1(141) <= to_unsigned(16#89#, 8);
  gmul3_1(142) <= to_unsigned(16#8A#, 8);
  gmul3_1(143) <= to_unsigned(16#AB#, 8);
  gmul3_1(144) <= to_unsigned(16#A8#, 8);
  gmul3_1(145) <= to_unsigned(16#AD#, 8);
  gmul3_1(146) <= to_unsigned(16#AE#, 8);
  gmul3_1(147) <= to_unsigned(16#A7#, 8);
  gmul3_1(148) <= to_unsigned(16#A4#, 8);
  gmul3_1(149) <= to_unsigned(16#A1#, 8);
  gmul3_1(150) <= to_unsigned(16#A2#, 8);
  gmul3_1(151) <= to_unsigned(16#B3#, 8);
  gmul3_1(152) <= to_unsigned(16#B0#, 8);
  gmul3_1(153) <= to_unsigned(16#B5#, 8);
  gmul3_1(154) <= to_unsigned(16#B6#, 8);
  gmul3_1(155) <= to_unsigned(16#BF#, 8);
  gmul3_1(156) <= to_unsigned(16#BC#, 8);
  gmul3_1(157) <= to_unsigned(16#B9#, 8);
  gmul3_1(158) <= to_unsigned(16#BA#, 8);
  gmul3_1(159) <= to_unsigned(16#FB#, 8);
  gmul3_1(160) <= to_unsigned(16#F8#, 8);
  gmul3_1(161) <= to_unsigned(16#FD#, 8);
  gmul3_1(162) <= to_unsigned(16#FE#, 8);
  gmul3_1(163) <= to_unsigned(16#F7#, 8);
  gmul3_1(164) <= to_unsigned(16#F4#, 8);
  gmul3_1(165) <= to_unsigned(16#F1#, 8);
  gmul3_1(166) <= to_unsigned(16#F2#, 8);
  gmul3_1(167) <= to_unsigned(16#E3#, 8);
  gmul3_1(168) <= to_unsigned(16#E0#, 8);
  gmul3_1(169) <= to_unsigned(16#E5#, 8);
  gmul3_1(170) <= to_unsigned(16#E6#, 8);
  gmul3_1(171) <= to_unsigned(16#EF#, 8);
  gmul3_1(172) <= to_unsigned(16#EC#, 8);
  gmul3_1(173) <= to_unsigned(16#E9#, 8);
  gmul3_1(174) <= to_unsigned(16#EA#, 8);
  gmul3_1(175) <= to_unsigned(16#CB#, 8);
  gmul3_1(176) <= to_unsigned(16#C8#, 8);
  gmul3_1(177) <= to_unsigned(16#CD#, 8);
  gmul3_1(178) <= to_unsigned(16#CE#, 8);
  gmul3_1(179) <= to_unsigned(16#C7#, 8);
  gmul3_1(180) <= to_unsigned(16#C4#, 8);
  gmul3_1(181) <= to_unsigned(16#C1#, 8);
  gmul3_1(182) <= to_unsigned(16#C2#, 8);
  gmul3_1(183) <= to_unsigned(16#D3#, 8);
  gmul3_1(184) <= to_unsigned(16#D0#, 8);
  gmul3_1(185) <= to_unsigned(16#D5#, 8);
  gmul3_1(186) <= to_unsigned(16#D6#, 8);
  gmul3_1(187) <= to_unsigned(16#DF#, 8);
  gmul3_1(188) <= to_unsigned(16#DC#, 8);
  gmul3_1(189) <= to_unsigned(16#D9#, 8);
  gmul3_1(190) <= to_unsigned(16#DA#, 8);
  gmul3_1(191) <= to_unsigned(16#5B#, 8);
  gmul3_1(192) <= to_unsigned(16#58#, 8);
  gmul3_1(193) <= to_unsigned(16#5D#, 8);
  gmul3_1(194) <= to_unsigned(16#5E#, 8);
  gmul3_1(195) <= to_unsigned(16#57#, 8);
  gmul3_1(196) <= to_unsigned(16#54#, 8);
  gmul3_1(197) <= to_unsigned(16#51#, 8);
  gmul3_1(198) <= to_unsigned(16#52#, 8);
  gmul3_1(199) <= to_unsigned(16#43#, 8);
  gmul3_1(200) <= to_unsigned(16#40#, 8);
  gmul3_1(201) <= to_unsigned(16#45#, 8);
  gmul3_1(202) <= to_unsigned(16#46#, 8);
  gmul3_1(203) <= to_unsigned(16#4F#, 8);
  gmul3_1(204) <= to_unsigned(16#4C#, 8);
  gmul3_1(205) <= to_unsigned(16#49#, 8);
  gmul3_1(206) <= to_unsigned(16#4A#, 8);
  gmul3_1(207) <= to_unsigned(16#6B#, 8);
  gmul3_1(208) <= to_unsigned(16#68#, 8);
  gmul3_1(209) <= to_unsigned(16#6D#, 8);
  gmul3_1(210) <= to_unsigned(16#6E#, 8);
  gmul3_1(211) <= to_unsigned(16#67#, 8);
  gmul3_1(212) <= to_unsigned(16#64#, 8);
  gmul3_1(213) <= to_unsigned(16#61#, 8);
  gmul3_1(214) <= to_unsigned(16#62#, 8);
  gmul3_1(215) <= to_unsigned(16#73#, 8);
  gmul3_1(216) <= to_unsigned(16#70#, 8);
  gmul3_1(217) <= to_unsigned(16#75#, 8);
  gmul3_1(218) <= to_unsigned(16#76#, 8);
  gmul3_1(219) <= to_unsigned(16#7F#, 8);
  gmul3_1(220) <= to_unsigned(16#7C#, 8);
  gmul3_1(221) <= to_unsigned(16#79#, 8);
  gmul3_1(222) <= to_unsigned(16#7A#, 8);
  gmul3_1(223) <= to_unsigned(16#3B#, 8);
  gmul3_1(224) <= to_unsigned(16#38#, 8);
  gmul3_1(225) <= to_unsigned(16#3D#, 8);
  gmul3_1(226) <= to_unsigned(16#3E#, 8);
  gmul3_1(227) <= to_unsigned(16#37#, 8);
  gmul3_1(228) <= to_unsigned(16#34#, 8);
  gmul3_1(229) <= to_unsigned(16#31#, 8);
  gmul3_1(230) <= to_unsigned(16#32#, 8);
  gmul3_1(231) <= to_unsigned(16#23#, 8);
  gmul3_1(232) <= to_unsigned(16#20#, 8);
  gmul3_1(233) <= to_unsigned(16#25#, 8);
  gmul3_1(234) <= to_unsigned(16#26#, 8);
  gmul3_1(235) <= to_unsigned(16#2F#, 8);
  gmul3_1(236) <= to_unsigned(16#2C#, 8);
  gmul3_1(237) <= to_unsigned(16#29#, 8);
  gmul3_1(238) <= to_unsigned(16#2A#, 8);
  gmul3_1(239) <= to_unsigned(16#0B#, 8);
  gmul3_1(240) <= to_unsigned(16#08#, 8);
  gmul3_1(241) <= to_unsigned(16#0D#, 8);
  gmul3_1(242) <= to_unsigned(16#0E#, 8);
  gmul3_1(243) <= to_unsigned(16#07#, 8);
  gmul3_1(244) <= to_unsigned(16#04#, 8);
  gmul3_1(245) <= to_unsigned(16#01#, 8);
  gmul3_1(246) <= to_unsigned(16#02#, 8);
  gmul3_1(247) <= to_unsigned(16#13#, 8);
  gmul3_1(248) <= to_unsigned(16#10#, 8);
  gmul3_1(249) <= to_unsigned(16#15#, 8);
  gmul3_1(250) <= to_unsigned(16#16#, 8);
  gmul3_1(251) <= to_unsigned(16#1F#, 8);
  gmul3_1(252) <= to_unsigned(16#1C#, 8);
  gmul3_1(253) <= to_unsigned(16#19#, 8);
  gmul3_1(254) <= to_unsigned(16#1A#, 8);
  gmul3_1(255) <= to_unsigned(16#1A#, 8);

  gmul2_2(0) <= to_unsigned(16#02#, 8);
  gmul2_2(1) <= to_unsigned(16#04#, 8);
  gmul2_2(2) <= to_unsigned(16#06#, 8);
  gmul2_2(3) <= to_unsigned(16#08#, 8);
  gmul2_2(4) <= to_unsigned(16#0A#, 8);
  gmul2_2(5) <= to_unsigned(16#0C#, 8);
  gmul2_2(6) <= to_unsigned(16#0E#, 8);
  gmul2_2(7) <= to_unsigned(16#10#, 8);
  gmul2_2(8) <= to_unsigned(16#12#, 8);
  gmul2_2(9) <= to_unsigned(16#14#, 8);
  gmul2_2(10) <= to_unsigned(16#16#, 8);
  gmul2_2(11) <= to_unsigned(16#18#, 8);
  gmul2_2(12) <= to_unsigned(16#1A#, 8);
  gmul2_2(13) <= to_unsigned(16#1C#, 8);
  gmul2_2(14) <= to_unsigned(16#1E#, 8);
  gmul2_2(15) <= to_unsigned(16#20#, 8);
  gmul2_2(16) <= to_unsigned(16#22#, 8);
  gmul2_2(17) <= to_unsigned(16#24#, 8);
  gmul2_2(18) <= to_unsigned(16#26#, 8);
  gmul2_2(19) <= to_unsigned(16#28#, 8);
  gmul2_2(20) <= to_unsigned(16#2A#, 8);
  gmul2_2(21) <= to_unsigned(16#2C#, 8);
  gmul2_2(22) <= to_unsigned(16#2E#, 8);
  gmul2_2(23) <= to_unsigned(16#30#, 8);
  gmul2_2(24) <= to_unsigned(16#32#, 8);
  gmul2_2(25) <= to_unsigned(16#34#, 8);
  gmul2_2(26) <= to_unsigned(16#36#, 8);
  gmul2_2(27) <= to_unsigned(16#38#, 8);
  gmul2_2(28) <= to_unsigned(16#3A#, 8);
  gmul2_2(29) <= to_unsigned(16#3C#, 8);
  gmul2_2(30) <= to_unsigned(16#3E#, 8);
  gmul2_2(31) <= to_unsigned(16#40#, 8);
  gmul2_2(32) <= to_unsigned(16#42#, 8);
  gmul2_2(33) <= to_unsigned(16#44#, 8);
  gmul2_2(34) <= to_unsigned(16#46#, 8);
  gmul2_2(35) <= to_unsigned(16#48#, 8);
  gmul2_2(36) <= to_unsigned(16#4A#, 8);
  gmul2_2(37) <= to_unsigned(16#4C#, 8);
  gmul2_2(38) <= to_unsigned(16#4E#, 8);
  gmul2_2(39) <= to_unsigned(16#50#, 8);
  gmul2_2(40) <= to_unsigned(16#52#, 8);
  gmul2_2(41) <= to_unsigned(16#54#, 8);
  gmul2_2(42) <= to_unsigned(16#56#, 8);
  gmul2_2(43) <= to_unsigned(16#58#, 8);
  gmul2_2(44) <= to_unsigned(16#5A#, 8);
  gmul2_2(45) <= to_unsigned(16#5C#, 8);
  gmul2_2(46) <= to_unsigned(16#5E#, 8);
  gmul2_2(47) <= to_unsigned(16#60#, 8);
  gmul2_2(48) <= to_unsigned(16#62#, 8);
  gmul2_2(49) <= to_unsigned(16#64#, 8);
  gmul2_2(50) <= to_unsigned(16#66#, 8);
  gmul2_2(51) <= to_unsigned(16#68#, 8);
  gmul2_2(52) <= to_unsigned(16#6A#, 8);
  gmul2_2(53) <= to_unsigned(16#6C#, 8);
  gmul2_2(54) <= to_unsigned(16#6E#, 8);
  gmul2_2(55) <= to_unsigned(16#70#, 8);
  gmul2_2(56) <= to_unsigned(16#72#, 8);
  gmul2_2(57) <= to_unsigned(16#74#, 8);
  gmul2_2(58) <= to_unsigned(16#76#, 8);
  gmul2_2(59) <= to_unsigned(16#78#, 8);
  gmul2_2(60) <= to_unsigned(16#7A#, 8);
  gmul2_2(61) <= to_unsigned(16#7C#, 8);
  gmul2_2(62) <= to_unsigned(16#7E#, 8);
  gmul2_2(63) <= to_unsigned(16#80#, 8);
  gmul2_2(64) <= to_unsigned(16#82#, 8);
  gmul2_2(65) <= to_unsigned(16#84#, 8);
  gmul2_2(66) <= to_unsigned(16#86#, 8);
  gmul2_2(67) <= to_unsigned(16#88#, 8);
  gmul2_2(68) <= to_unsigned(16#8A#, 8);
  gmul2_2(69) <= to_unsigned(16#8C#, 8);
  gmul2_2(70) <= to_unsigned(16#8E#, 8);
  gmul2_2(71) <= to_unsigned(16#90#, 8);
  gmul2_2(72) <= to_unsigned(16#92#, 8);
  gmul2_2(73) <= to_unsigned(16#94#, 8);
  gmul2_2(74) <= to_unsigned(16#96#, 8);
  gmul2_2(75) <= to_unsigned(16#98#, 8);
  gmul2_2(76) <= to_unsigned(16#9A#, 8);
  gmul2_2(77) <= to_unsigned(16#9C#, 8);
  gmul2_2(78) <= to_unsigned(16#9E#, 8);
  gmul2_2(79) <= to_unsigned(16#A0#, 8);
  gmul2_2(80) <= to_unsigned(16#A2#, 8);
  gmul2_2(81) <= to_unsigned(16#A4#, 8);
  gmul2_2(82) <= to_unsigned(16#A6#, 8);
  gmul2_2(83) <= to_unsigned(16#A8#, 8);
  gmul2_2(84) <= to_unsigned(16#AA#, 8);
  gmul2_2(85) <= to_unsigned(16#AC#, 8);
  gmul2_2(86) <= to_unsigned(16#AE#, 8);
  gmul2_2(87) <= to_unsigned(16#B0#, 8);
  gmul2_2(88) <= to_unsigned(16#B2#, 8);
  gmul2_2(89) <= to_unsigned(16#B4#, 8);
  gmul2_2(90) <= to_unsigned(16#B6#, 8);
  gmul2_2(91) <= to_unsigned(16#B8#, 8);
  gmul2_2(92) <= to_unsigned(16#BA#, 8);
  gmul2_2(93) <= to_unsigned(16#BC#, 8);
  gmul2_2(94) <= to_unsigned(16#BE#, 8);
  gmul2_2(95) <= to_unsigned(16#C0#, 8);
  gmul2_2(96) <= to_unsigned(16#C2#, 8);
  gmul2_2(97) <= to_unsigned(16#C4#, 8);
  gmul2_2(98) <= to_unsigned(16#C6#, 8);
  gmul2_2(99) <= to_unsigned(16#C8#, 8);
  gmul2_2(100) <= to_unsigned(16#CA#, 8);
  gmul2_2(101) <= to_unsigned(16#CC#, 8);
  gmul2_2(102) <= to_unsigned(16#CE#, 8);
  gmul2_2(103) <= to_unsigned(16#D0#, 8);
  gmul2_2(104) <= to_unsigned(16#D2#, 8);
  gmul2_2(105) <= to_unsigned(16#D4#, 8);
  gmul2_2(106) <= to_unsigned(16#D6#, 8);
  gmul2_2(107) <= to_unsigned(16#D8#, 8);
  gmul2_2(108) <= to_unsigned(16#DA#, 8);
  gmul2_2(109) <= to_unsigned(16#DC#, 8);
  gmul2_2(110) <= to_unsigned(16#DE#, 8);
  gmul2_2(111) <= to_unsigned(16#E0#, 8);
  gmul2_2(112) <= to_unsigned(16#E2#, 8);
  gmul2_2(113) <= to_unsigned(16#E4#, 8);
  gmul2_2(114) <= to_unsigned(16#E6#, 8);
  gmul2_2(115) <= to_unsigned(16#E8#, 8);
  gmul2_2(116) <= to_unsigned(16#EA#, 8);
  gmul2_2(117) <= to_unsigned(16#EC#, 8);
  gmul2_2(118) <= to_unsigned(16#EE#, 8);
  gmul2_2(119) <= to_unsigned(16#F0#, 8);
  gmul2_2(120) <= to_unsigned(16#F2#, 8);
  gmul2_2(121) <= to_unsigned(16#F4#, 8);
  gmul2_2(122) <= to_unsigned(16#F6#, 8);
  gmul2_2(123) <= to_unsigned(16#F8#, 8);
  gmul2_2(124) <= to_unsigned(16#FA#, 8);
  gmul2_2(125) <= to_unsigned(16#FC#, 8);
  gmul2_2(126) <= to_unsigned(16#FE#, 8);
  gmul2_2(127) <= to_unsigned(16#1B#, 8);
  gmul2_2(128) <= to_unsigned(16#19#, 8);
  gmul2_2(129) <= to_unsigned(16#1F#, 8);
  gmul2_2(130) <= to_unsigned(16#1D#, 8);
  gmul2_2(131) <= to_unsigned(16#13#, 8);
  gmul2_2(132) <= to_unsigned(16#11#, 8);
  gmul2_2(133) <= to_unsigned(16#17#, 8);
  gmul2_2(134) <= to_unsigned(16#15#, 8);
  gmul2_2(135) <= to_unsigned(16#0B#, 8);
  gmul2_2(136) <= to_unsigned(16#09#, 8);
  gmul2_2(137) <= to_unsigned(16#0F#, 8);
  gmul2_2(138) <= to_unsigned(16#0D#, 8);
  gmul2_2(139) <= to_unsigned(16#03#, 8);
  gmul2_2(140) <= to_unsigned(16#01#, 8);
  gmul2_2(141) <= to_unsigned(16#07#, 8);
  gmul2_2(142) <= to_unsigned(16#05#, 8);
  gmul2_2(143) <= to_unsigned(16#3B#, 8);
  gmul2_2(144) <= to_unsigned(16#39#, 8);
  gmul2_2(145) <= to_unsigned(16#3F#, 8);
  gmul2_2(146) <= to_unsigned(16#3D#, 8);
  gmul2_2(147) <= to_unsigned(16#33#, 8);
  gmul2_2(148) <= to_unsigned(16#31#, 8);
  gmul2_2(149) <= to_unsigned(16#37#, 8);
  gmul2_2(150) <= to_unsigned(16#35#, 8);
  gmul2_2(151) <= to_unsigned(16#2B#, 8);
  gmul2_2(152) <= to_unsigned(16#29#, 8);
  gmul2_2(153) <= to_unsigned(16#2F#, 8);
  gmul2_2(154) <= to_unsigned(16#2D#, 8);
  gmul2_2(155) <= to_unsigned(16#23#, 8);
  gmul2_2(156) <= to_unsigned(16#21#, 8);
  gmul2_2(157) <= to_unsigned(16#27#, 8);
  gmul2_2(158) <= to_unsigned(16#25#, 8);
  gmul2_2(159) <= to_unsigned(16#5B#, 8);
  gmul2_2(160) <= to_unsigned(16#59#, 8);
  gmul2_2(161) <= to_unsigned(16#5F#, 8);
  gmul2_2(162) <= to_unsigned(16#5D#, 8);
  gmul2_2(163) <= to_unsigned(16#53#, 8);
  gmul2_2(164) <= to_unsigned(16#51#, 8);
  gmul2_2(165) <= to_unsigned(16#57#, 8);
  gmul2_2(166) <= to_unsigned(16#55#, 8);
  gmul2_2(167) <= to_unsigned(16#4B#, 8);
  gmul2_2(168) <= to_unsigned(16#49#, 8);
  gmul2_2(169) <= to_unsigned(16#4F#, 8);
  gmul2_2(170) <= to_unsigned(16#4D#, 8);
  gmul2_2(171) <= to_unsigned(16#43#, 8);
  gmul2_2(172) <= to_unsigned(16#41#, 8);
  gmul2_2(173) <= to_unsigned(16#47#, 8);
  gmul2_2(174) <= to_unsigned(16#45#, 8);
  gmul2_2(175) <= to_unsigned(16#7B#, 8);
  gmul2_2(176) <= to_unsigned(16#79#, 8);
  gmul2_2(177) <= to_unsigned(16#7F#, 8);
  gmul2_2(178) <= to_unsigned(16#7D#, 8);
  gmul2_2(179) <= to_unsigned(16#73#, 8);
  gmul2_2(180) <= to_unsigned(16#71#, 8);
  gmul2_2(181) <= to_unsigned(16#77#, 8);
  gmul2_2(182) <= to_unsigned(16#75#, 8);
  gmul2_2(183) <= to_unsigned(16#6B#, 8);
  gmul2_2(184) <= to_unsigned(16#69#, 8);
  gmul2_2(185) <= to_unsigned(16#6F#, 8);
  gmul2_2(186) <= to_unsigned(16#6D#, 8);
  gmul2_2(187) <= to_unsigned(16#63#, 8);
  gmul2_2(188) <= to_unsigned(16#61#, 8);
  gmul2_2(189) <= to_unsigned(16#67#, 8);
  gmul2_2(190) <= to_unsigned(16#65#, 8);
  gmul2_2(191) <= to_unsigned(16#9B#, 8);
  gmul2_2(192) <= to_unsigned(16#99#, 8);
  gmul2_2(193) <= to_unsigned(16#9F#, 8);
  gmul2_2(194) <= to_unsigned(16#9D#, 8);
  gmul2_2(195) <= to_unsigned(16#93#, 8);
  gmul2_2(196) <= to_unsigned(16#91#, 8);
  gmul2_2(197) <= to_unsigned(16#97#, 8);
  gmul2_2(198) <= to_unsigned(16#95#, 8);
  gmul2_2(199) <= to_unsigned(16#8B#, 8);
  gmul2_2(200) <= to_unsigned(16#89#, 8);
  gmul2_2(201) <= to_unsigned(16#8F#, 8);
  gmul2_2(202) <= to_unsigned(16#8D#, 8);
  gmul2_2(203) <= to_unsigned(16#83#, 8);
  gmul2_2(204) <= to_unsigned(16#81#, 8);
  gmul2_2(205) <= to_unsigned(16#87#, 8);
  gmul2_2(206) <= to_unsigned(16#85#, 8);
  gmul2_2(207) <= to_unsigned(16#BB#, 8);
  gmul2_2(208) <= to_unsigned(16#B9#, 8);
  gmul2_2(209) <= to_unsigned(16#BF#, 8);
  gmul2_2(210) <= to_unsigned(16#BD#, 8);
  gmul2_2(211) <= to_unsigned(16#B3#, 8);
  gmul2_2(212) <= to_unsigned(16#B1#, 8);
  gmul2_2(213) <= to_unsigned(16#B7#, 8);
  gmul2_2(214) <= to_unsigned(16#B5#, 8);
  gmul2_2(215) <= to_unsigned(16#AB#, 8);
  gmul2_2(216) <= to_unsigned(16#A9#, 8);
  gmul2_2(217) <= to_unsigned(16#AF#, 8);
  gmul2_2(218) <= to_unsigned(16#AD#, 8);
  gmul2_2(219) <= to_unsigned(16#A3#, 8);
  gmul2_2(220) <= to_unsigned(16#A1#, 8);
  gmul2_2(221) <= to_unsigned(16#A7#, 8);
  gmul2_2(222) <= to_unsigned(16#A5#, 8);
  gmul2_2(223) <= to_unsigned(16#DB#, 8);
  gmul2_2(224) <= to_unsigned(16#D9#, 8);
  gmul2_2(225) <= to_unsigned(16#DF#, 8);
  gmul2_2(226) <= to_unsigned(16#DD#, 8);
  gmul2_2(227) <= to_unsigned(16#D3#, 8);
  gmul2_2(228) <= to_unsigned(16#D1#, 8);
  gmul2_2(229) <= to_unsigned(16#D7#, 8);
  gmul2_2(230) <= to_unsigned(16#D5#, 8);
  gmul2_2(231) <= to_unsigned(16#CB#, 8);
  gmul2_2(232) <= to_unsigned(16#C9#, 8);
  gmul2_2(233) <= to_unsigned(16#CF#, 8);
  gmul2_2(234) <= to_unsigned(16#CD#, 8);
  gmul2_2(235) <= to_unsigned(16#C3#, 8);
  gmul2_2(236) <= to_unsigned(16#C1#, 8);
  gmul2_2(237) <= to_unsigned(16#C7#, 8);
  gmul2_2(238) <= to_unsigned(16#C5#, 8);
  gmul2_2(239) <= to_unsigned(16#FB#, 8);
  gmul2_2(240) <= to_unsigned(16#F9#, 8);
  gmul2_2(241) <= to_unsigned(16#FF#, 8);
  gmul2_2(242) <= to_unsigned(16#FD#, 8);
  gmul2_2(243) <= to_unsigned(16#F3#, 8);
  gmul2_2(244) <= to_unsigned(16#F1#, 8);
  gmul2_2(245) <= to_unsigned(16#F7#, 8);
  gmul2_2(246) <= to_unsigned(16#F5#, 8);
  gmul2_2(247) <= to_unsigned(16#EB#, 8);
  gmul2_2(248) <= to_unsigned(16#E9#, 8);
  gmul2_2(249) <= to_unsigned(16#EF#, 8);
  gmul2_2(250) <= to_unsigned(16#ED#, 8);
  gmul2_2(251) <= to_unsigned(16#E3#, 8);
  gmul2_2(252) <= to_unsigned(16#E1#, 8);
  gmul2_2(253) <= to_unsigned(16#E7#, 8);
  gmul2_2(254) <= to_unsigned(16#E5#, 8);
  gmul2_2(255) <= to_unsigned(16#E5#, 8);

  gmul3_2(0) <= to_unsigned(16#03#, 8);
  gmul3_2(1) <= to_unsigned(16#06#, 8);
  gmul3_2(2) <= to_unsigned(16#05#, 8);
  gmul3_2(3) <= to_unsigned(16#0C#, 8);
  gmul3_2(4) <= to_unsigned(16#0F#, 8);
  gmul3_2(5) <= to_unsigned(16#0A#, 8);
  gmul3_2(6) <= to_unsigned(16#09#, 8);
  gmul3_2(7) <= to_unsigned(16#18#, 8);
  gmul3_2(8) <= to_unsigned(16#1B#, 8);
  gmul3_2(9) <= to_unsigned(16#1E#, 8);
  gmul3_2(10) <= to_unsigned(16#1D#, 8);
  gmul3_2(11) <= to_unsigned(16#14#, 8);
  gmul3_2(12) <= to_unsigned(16#17#, 8);
  gmul3_2(13) <= to_unsigned(16#12#, 8);
  gmul3_2(14) <= to_unsigned(16#11#, 8);
  gmul3_2(15) <= to_unsigned(16#30#, 8);
  gmul3_2(16) <= to_unsigned(16#33#, 8);
  gmul3_2(17) <= to_unsigned(16#36#, 8);
  gmul3_2(18) <= to_unsigned(16#35#, 8);
  gmul3_2(19) <= to_unsigned(16#3C#, 8);
  gmul3_2(20) <= to_unsigned(16#3F#, 8);
  gmul3_2(21) <= to_unsigned(16#3A#, 8);
  gmul3_2(22) <= to_unsigned(16#39#, 8);
  gmul3_2(23) <= to_unsigned(16#28#, 8);
  gmul3_2(24) <= to_unsigned(16#2B#, 8);
  gmul3_2(25) <= to_unsigned(16#2E#, 8);
  gmul3_2(26) <= to_unsigned(16#2D#, 8);
  gmul3_2(27) <= to_unsigned(16#24#, 8);
  gmul3_2(28) <= to_unsigned(16#27#, 8);
  gmul3_2(29) <= to_unsigned(16#22#, 8);
  gmul3_2(30) <= to_unsigned(16#21#, 8);
  gmul3_2(31) <= to_unsigned(16#60#, 8);
  gmul3_2(32) <= to_unsigned(16#63#, 8);
  gmul3_2(33) <= to_unsigned(16#66#, 8);
  gmul3_2(34) <= to_unsigned(16#65#, 8);
  gmul3_2(35) <= to_unsigned(16#6C#, 8);
  gmul3_2(36) <= to_unsigned(16#6F#, 8);
  gmul3_2(37) <= to_unsigned(16#6A#, 8);
  gmul3_2(38) <= to_unsigned(16#69#, 8);
  gmul3_2(39) <= to_unsigned(16#78#, 8);
  gmul3_2(40) <= to_unsigned(16#7B#, 8);
  gmul3_2(41) <= to_unsigned(16#7E#, 8);
  gmul3_2(42) <= to_unsigned(16#7D#, 8);
  gmul3_2(43) <= to_unsigned(16#74#, 8);
  gmul3_2(44) <= to_unsigned(16#77#, 8);
  gmul3_2(45) <= to_unsigned(16#72#, 8);
  gmul3_2(46) <= to_unsigned(16#71#, 8);
  gmul3_2(47) <= to_unsigned(16#50#, 8);
  gmul3_2(48) <= to_unsigned(16#53#, 8);
  gmul3_2(49) <= to_unsigned(16#56#, 8);
  gmul3_2(50) <= to_unsigned(16#55#, 8);
  gmul3_2(51) <= to_unsigned(16#5C#, 8);
  gmul3_2(52) <= to_unsigned(16#5F#, 8);
  gmul3_2(53) <= to_unsigned(16#5A#, 8);
  gmul3_2(54) <= to_unsigned(16#59#, 8);
  gmul3_2(55) <= to_unsigned(16#48#, 8);
  gmul3_2(56) <= to_unsigned(16#4B#, 8);
  gmul3_2(57) <= to_unsigned(16#4E#, 8);
  gmul3_2(58) <= to_unsigned(16#4D#, 8);
  gmul3_2(59) <= to_unsigned(16#44#, 8);
  gmul3_2(60) <= to_unsigned(16#47#, 8);
  gmul3_2(61) <= to_unsigned(16#42#, 8);
  gmul3_2(62) <= to_unsigned(16#41#, 8);
  gmul3_2(63) <= to_unsigned(16#C0#, 8);
  gmul3_2(64) <= to_unsigned(16#C3#, 8);
  gmul3_2(65) <= to_unsigned(16#C6#, 8);
  gmul3_2(66) <= to_unsigned(16#C5#, 8);
  gmul3_2(67) <= to_unsigned(16#CC#, 8);
  gmul3_2(68) <= to_unsigned(16#CF#, 8);
  gmul3_2(69) <= to_unsigned(16#CA#, 8);
  gmul3_2(70) <= to_unsigned(16#C9#, 8);
  gmul3_2(71) <= to_unsigned(16#D8#, 8);
  gmul3_2(72) <= to_unsigned(16#DB#, 8);
  gmul3_2(73) <= to_unsigned(16#DE#, 8);
  gmul3_2(74) <= to_unsigned(16#DD#, 8);
  gmul3_2(75) <= to_unsigned(16#D4#, 8);
  gmul3_2(76) <= to_unsigned(16#D7#, 8);
  gmul3_2(77) <= to_unsigned(16#D2#, 8);
  gmul3_2(78) <= to_unsigned(16#D1#, 8);
  gmul3_2(79) <= to_unsigned(16#F0#, 8);
  gmul3_2(80) <= to_unsigned(16#F3#, 8);
  gmul3_2(81) <= to_unsigned(16#F6#, 8);
  gmul3_2(82) <= to_unsigned(16#F5#, 8);
  gmul3_2(83) <= to_unsigned(16#FC#, 8);
  gmul3_2(84) <= to_unsigned(16#FF#, 8);
  gmul3_2(85) <= to_unsigned(16#FA#, 8);
  gmul3_2(86) <= to_unsigned(16#F9#, 8);
  gmul3_2(87) <= to_unsigned(16#E8#, 8);
  gmul3_2(88) <= to_unsigned(16#EB#, 8);
  gmul3_2(89) <= to_unsigned(16#EE#, 8);
  gmul3_2(90) <= to_unsigned(16#ED#, 8);
  gmul3_2(91) <= to_unsigned(16#E4#, 8);
  gmul3_2(92) <= to_unsigned(16#E7#, 8);
  gmul3_2(93) <= to_unsigned(16#E2#, 8);
  gmul3_2(94) <= to_unsigned(16#E1#, 8);
  gmul3_2(95) <= to_unsigned(16#A0#, 8);
  gmul3_2(96) <= to_unsigned(16#A3#, 8);
  gmul3_2(97) <= to_unsigned(16#A6#, 8);
  gmul3_2(98) <= to_unsigned(16#A5#, 8);
  gmul3_2(99) <= to_unsigned(16#AC#, 8);
  gmul3_2(100) <= to_unsigned(16#AF#, 8);
  gmul3_2(101) <= to_unsigned(16#AA#, 8);
  gmul3_2(102) <= to_unsigned(16#A9#, 8);
  gmul3_2(103) <= to_unsigned(16#B8#, 8);
  gmul3_2(104) <= to_unsigned(16#BB#, 8);
  gmul3_2(105) <= to_unsigned(16#BE#, 8);
  gmul3_2(106) <= to_unsigned(16#BD#, 8);
  gmul3_2(107) <= to_unsigned(16#B4#, 8);
  gmul3_2(108) <= to_unsigned(16#B7#, 8);
  gmul3_2(109) <= to_unsigned(16#B2#, 8);
  gmul3_2(110) <= to_unsigned(16#B1#, 8);
  gmul3_2(111) <= to_unsigned(16#90#, 8);
  gmul3_2(112) <= to_unsigned(16#93#, 8);
  gmul3_2(113) <= to_unsigned(16#96#, 8);
  gmul3_2(114) <= to_unsigned(16#95#, 8);
  gmul3_2(115) <= to_unsigned(16#9C#, 8);
  gmul3_2(116) <= to_unsigned(16#9F#, 8);
  gmul3_2(117) <= to_unsigned(16#9A#, 8);
  gmul3_2(118) <= to_unsigned(16#99#, 8);
  gmul3_2(119) <= to_unsigned(16#88#, 8);
  gmul3_2(120) <= to_unsigned(16#8B#, 8);
  gmul3_2(121) <= to_unsigned(16#8E#, 8);
  gmul3_2(122) <= to_unsigned(16#8D#, 8);
  gmul3_2(123) <= to_unsigned(16#84#, 8);
  gmul3_2(124) <= to_unsigned(16#87#, 8);
  gmul3_2(125) <= to_unsigned(16#82#, 8);
  gmul3_2(126) <= to_unsigned(16#81#, 8);
  gmul3_2(127) <= to_unsigned(16#9B#, 8);
  gmul3_2(128) <= to_unsigned(16#98#, 8);
  gmul3_2(129) <= to_unsigned(16#9D#, 8);
  gmul3_2(130) <= to_unsigned(16#9E#, 8);
  gmul3_2(131) <= to_unsigned(16#97#, 8);
  gmul3_2(132) <= to_unsigned(16#94#, 8);
  gmul3_2(133) <= to_unsigned(16#91#, 8);
  gmul3_2(134) <= to_unsigned(16#92#, 8);
  gmul3_2(135) <= to_unsigned(16#83#, 8);
  gmul3_2(136) <= to_unsigned(16#80#, 8);
  gmul3_2(137) <= to_unsigned(16#85#, 8);
  gmul3_2(138) <= to_unsigned(16#86#, 8);
  gmul3_2(139) <= to_unsigned(16#8F#, 8);
  gmul3_2(140) <= to_unsigned(16#8C#, 8);
  gmul3_2(141) <= to_unsigned(16#89#, 8);
  gmul3_2(142) <= to_unsigned(16#8A#, 8);
  gmul3_2(143) <= to_unsigned(16#AB#, 8);
  gmul3_2(144) <= to_unsigned(16#A8#, 8);
  gmul3_2(145) <= to_unsigned(16#AD#, 8);
  gmul3_2(146) <= to_unsigned(16#AE#, 8);
  gmul3_2(147) <= to_unsigned(16#A7#, 8);
  gmul3_2(148) <= to_unsigned(16#A4#, 8);
  gmul3_2(149) <= to_unsigned(16#A1#, 8);
  gmul3_2(150) <= to_unsigned(16#A2#, 8);
  gmul3_2(151) <= to_unsigned(16#B3#, 8);
  gmul3_2(152) <= to_unsigned(16#B0#, 8);
  gmul3_2(153) <= to_unsigned(16#B5#, 8);
  gmul3_2(154) <= to_unsigned(16#B6#, 8);
  gmul3_2(155) <= to_unsigned(16#BF#, 8);
  gmul3_2(156) <= to_unsigned(16#BC#, 8);
  gmul3_2(157) <= to_unsigned(16#B9#, 8);
  gmul3_2(158) <= to_unsigned(16#BA#, 8);
  gmul3_2(159) <= to_unsigned(16#FB#, 8);
  gmul3_2(160) <= to_unsigned(16#F8#, 8);
  gmul3_2(161) <= to_unsigned(16#FD#, 8);
  gmul3_2(162) <= to_unsigned(16#FE#, 8);
  gmul3_2(163) <= to_unsigned(16#F7#, 8);
  gmul3_2(164) <= to_unsigned(16#F4#, 8);
  gmul3_2(165) <= to_unsigned(16#F1#, 8);
  gmul3_2(166) <= to_unsigned(16#F2#, 8);
  gmul3_2(167) <= to_unsigned(16#E3#, 8);
  gmul3_2(168) <= to_unsigned(16#E0#, 8);
  gmul3_2(169) <= to_unsigned(16#E5#, 8);
  gmul3_2(170) <= to_unsigned(16#E6#, 8);
  gmul3_2(171) <= to_unsigned(16#EF#, 8);
  gmul3_2(172) <= to_unsigned(16#EC#, 8);
  gmul3_2(173) <= to_unsigned(16#E9#, 8);
  gmul3_2(174) <= to_unsigned(16#EA#, 8);
  gmul3_2(175) <= to_unsigned(16#CB#, 8);
  gmul3_2(176) <= to_unsigned(16#C8#, 8);
  gmul3_2(177) <= to_unsigned(16#CD#, 8);
  gmul3_2(178) <= to_unsigned(16#CE#, 8);
  gmul3_2(179) <= to_unsigned(16#C7#, 8);
  gmul3_2(180) <= to_unsigned(16#C4#, 8);
  gmul3_2(181) <= to_unsigned(16#C1#, 8);
  gmul3_2(182) <= to_unsigned(16#C2#, 8);
  gmul3_2(183) <= to_unsigned(16#D3#, 8);
  gmul3_2(184) <= to_unsigned(16#D0#, 8);
  gmul3_2(185) <= to_unsigned(16#D5#, 8);
  gmul3_2(186) <= to_unsigned(16#D6#, 8);
  gmul3_2(187) <= to_unsigned(16#DF#, 8);
  gmul3_2(188) <= to_unsigned(16#DC#, 8);
  gmul3_2(189) <= to_unsigned(16#D9#, 8);
  gmul3_2(190) <= to_unsigned(16#DA#, 8);
  gmul3_2(191) <= to_unsigned(16#5B#, 8);
  gmul3_2(192) <= to_unsigned(16#58#, 8);
  gmul3_2(193) <= to_unsigned(16#5D#, 8);
  gmul3_2(194) <= to_unsigned(16#5E#, 8);
  gmul3_2(195) <= to_unsigned(16#57#, 8);
  gmul3_2(196) <= to_unsigned(16#54#, 8);
  gmul3_2(197) <= to_unsigned(16#51#, 8);
  gmul3_2(198) <= to_unsigned(16#52#, 8);
  gmul3_2(199) <= to_unsigned(16#43#, 8);
  gmul3_2(200) <= to_unsigned(16#40#, 8);
  gmul3_2(201) <= to_unsigned(16#45#, 8);
  gmul3_2(202) <= to_unsigned(16#46#, 8);
  gmul3_2(203) <= to_unsigned(16#4F#, 8);
  gmul3_2(204) <= to_unsigned(16#4C#, 8);
  gmul3_2(205) <= to_unsigned(16#49#, 8);
  gmul3_2(206) <= to_unsigned(16#4A#, 8);
  gmul3_2(207) <= to_unsigned(16#6B#, 8);
  gmul3_2(208) <= to_unsigned(16#68#, 8);
  gmul3_2(209) <= to_unsigned(16#6D#, 8);
  gmul3_2(210) <= to_unsigned(16#6E#, 8);
  gmul3_2(211) <= to_unsigned(16#67#, 8);
  gmul3_2(212) <= to_unsigned(16#64#, 8);
  gmul3_2(213) <= to_unsigned(16#61#, 8);
  gmul3_2(214) <= to_unsigned(16#62#, 8);
  gmul3_2(215) <= to_unsigned(16#73#, 8);
  gmul3_2(216) <= to_unsigned(16#70#, 8);
  gmul3_2(217) <= to_unsigned(16#75#, 8);
  gmul3_2(218) <= to_unsigned(16#76#, 8);
  gmul3_2(219) <= to_unsigned(16#7F#, 8);
  gmul3_2(220) <= to_unsigned(16#7C#, 8);
  gmul3_2(221) <= to_unsigned(16#79#, 8);
  gmul3_2(222) <= to_unsigned(16#7A#, 8);
  gmul3_2(223) <= to_unsigned(16#3B#, 8);
  gmul3_2(224) <= to_unsigned(16#38#, 8);
  gmul3_2(225) <= to_unsigned(16#3D#, 8);
  gmul3_2(226) <= to_unsigned(16#3E#, 8);
  gmul3_2(227) <= to_unsigned(16#37#, 8);
  gmul3_2(228) <= to_unsigned(16#34#, 8);
  gmul3_2(229) <= to_unsigned(16#31#, 8);
  gmul3_2(230) <= to_unsigned(16#32#, 8);
  gmul3_2(231) <= to_unsigned(16#23#, 8);
  gmul3_2(232) <= to_unsigned(16#20#, 8);
  gmul3_2(233) <= to_unsigned(16#25#, 8);
  gmul3_2(234) <= to_unsigned(16#26#, 8);
  gmul3_2(235) <= to_unsigned(16#2F#, 8);
  gmul3_2(236) <= to_unsigned(16#2C#, 8);
  gmul3_2(237) <= to_unsigned(16#29#, 8);
  gmul3_2(238) <= to_unsigned(16#2A#, 8);
  gmul3_2(239) <= to_unsigned(16#0B#, 8);
  gmul3_2(240) <= to_unsigned(16#08#, 8);
  gmul3_2(241) <= to_unsigned(16#0D#, 8);
  gmul3_2(242) <= to_unsigned(16#0E#, 8);
  gmul3_2(243) <= to_unsigned(16#07#, 8);
  gmul3_2(244) <= to_unsigned(16#04#, 8);
  gmul3_2(245) <= to_unsigned(16#01#, 8);
  gmul3_2(246) <= to_unsigned(16#02#, 8);
  gmul3_2(247) <= to_unsigned(16#13#, 8);
  gmul3_2(248) <= to_unsigned(16#10#, 8);
  gmul3_2(249) <= to_unsigned(16#15#, 8);
  gmul3_2(250) <= to_unsigned(16#16#, 8);
  gmul3_2(251) <= to_unsigned(16#1F#, 8);
  gmul3_2(252) <= to_unsigned(16#1C#, 8);
  gmul3_2(253) <= to_unsigned(16#19#, 8);
  gmul3_2(254) <= to_unsigned(16#1A#, 8);
  gmul3_2(255) <= to_unsigned(16#1A#, 8);

  gmul3_3(0) <= to_unsigned(16#03#, 8);
  gmul3_3(1) <= to_unsigned(16#06#, 8);
  gmul3_3(2) <= to_unsigned(16#05#, 8);
  gmul3_3(3) <= to_unsigned(16#0C#, 8);
  gmul3_3(4) <= to_unsigned(16#0F#, 8);
  gmul3_3(5) <= to_unsigned(16#0A#, 8);
  gmul3_3(6) <= to_unsigned(16#09#, 8);
  gmul3_3(7) <= to_unsigned(16#18#, 8);
  gmul3_3(8) <= to_unsigned(16#1B#, 8);
  gmul3_3(9) <= to_unsigned(16#1E#, 8);
  gmul3_3(10) <= to_unsigned(16#1D#, 8);
  gmul3_3(11) <= to_unsigned(16#14#, 8);
  gmul3_3(12) <= to_unsigned(16#17#, 8);
  gmul3_3(13) <= to_unsigned(16#12#, 8);
  gmul3_3(14) <= to_unsigned(16#11#, 8);
  gmul3_3(15) <= to_unsigned(16#30#, 8);
  gmul3_3(16) <= to_unsigned(16#33#, 8);
  gmul3_3(17) <= to_unsigned(16#36#, 8);
  gmul3_3(18) <= to_unsigned(16#35#, 8);
  gmul3_3(19) <= to_unsigned(16#3C#, 8);
  gmul3_3(20) <= to_unsigned(16#3F#, 8);
  gmul3_3(21) <= to_unsigned(16#3A#, 8);
  gmul3_3(22) <= to_unsigned(16#39#, 8);
  gmul3_3(23) <= to_unsigned(16#28#, 8);
  gmul3_3(24) <= to_unsigned(16#2B#, 8);
  gmul3_3(25) <= to_unsigned(16#2E#, 8);
  gmul3_3(26) <= to_unsigned(16#2D#, 8);
  gmul3_3(27) <= to_unsigned(16#24#, 8);
  gmul3_3(28) <= to_unsigned(16#27#, 8);
  gmul3_3(29) <= to_unsigned(16#22#, 8);
  gmul3_3(30) <= to_unsigned(16#21#, 8);
  gmul3_3(31) <= to_unsigned(16#60#, 8);
  gmul3_3(32) <= to_unsigned(16#63#, 8);
  gmul3_3(33) <= to_unsigned(16#66#, 8);
  gmul3_3(34) <= to_unsigned(16#65#, 8);
  gmul3_3(35) <= to_unsigned(16#6C#, 8);
  gmul3_3(36) <= to_unsigned(16#6F#, 8);
  gmul3_3(37) <= to_unsigned(16#6A#, 8);
  gmul3_3(38) <= to_unsigned(16#69#, 8);
  gmul3_3(39) <= to_unsigned(16#78#, 8);
  gmul3_3(40) <= to_unsigned(16#7B#, 8);
  gmul3_3(41) <= to_unsigned(16#7E#, 8);
  gmul3_3(42) <= to_unsigned(16#7D#, 8);
  gmul3_3(43) <= to_unsigned(16#74#, 8);
  gmul3_3(44) <= to_unsigned(16#77#, 8);
  gmul3_3(45) <= to_unsigned(16#72#, 8);
  gmul3_3(46) <= to_unsigned(16#71#, 8);
  gmul3_3(47) <= to_unsigned(16#50#, 8);
  gmul3_3(48) <= to_unsigned(16#53#, 8);
  gmul3_3(49) <= to_unsigned(16#56#, 8);
  gmul3_3(50) <= to_unsigned(16#55#, 8);
  gmul3_3(51) <= to_unsigned(16#5C#, 8);
  gmul3_3(52) <= to_unsigned(16#5F#, 8);
  gmul3_3(53) <= to_unsigned(16#5A#, 8);
  gmul3_3(54) <= to_unsigned(16#59#, 8);
  gmul3_3(55) <= to_unsigned(16#48#, 8);
  gmul3_3(56) <= to_unsigned(16#4B#, 8);
  gmul3_3(57) <= to_unsigned(16#4E#, 8);
  gmul3_3(58) <= to_unsigned(16#4D#, 8);
  gmul3_3(59) <= to_unsigned(16#44#, 8);
  gmul3_3(60) <= to_unsigned(16#47#, 8);
  gmul3_3(61) <= to_unsigned(16#42#, 8);
  gmul3_3(62) <= to_unsigned(16#41#, 8);
  gmul3_3(63) <= to_unsigned(16#C0#, 8);
  gmul3_3(64) <= to_unsigned(16#C3#, 8);
  gmul3_3(65) <= to_unsigned(16#C6#, 8);
  gmul3_3(66) <= to_unsigned(16#C5#, 8);
  gmul3_3(67) <= to_unsigned(16#CC#, 8);
  gmul3_3(68) <= to_unsigned(16#CF#, 8);
  gmul3_3(69) <= to_unsigned(16#CA#, 8);
  gmul3_3(70) <= to_unsigned(16#C9#, 8);
  gmul3_3(71) <= to_unsigned(16#D8#, 8);
  gmul3_3(72) <= to_unsigned(16#DB#, 8);
  gmul3_3(73) <= to_unsigned(16#DE#, 8);
  gmul3_3(74) <= to_unsigned(16#DD#, 8);
  gmul3_3(75) <= to_unsigned(16#D4#, 8);
  gmul3_3(76) <= to_unsigned(16#D7#, 8);
  gmul3_3(77) <= to_unsigned(16#D2#, 8);
  gmul3_3(78) <= to_unsigned(16#D1#, 8);
  gmul3_3(79) <= to_unsigned(16#F0#, 8);
  gmul3_3(80) <= to_unsigned(16#F3#, 8);
  gmul3_3(81) <= to_unsigned(16#F6#, 8);
  gmul3_3(82) <= to_unsigned(16#F5#, 8);
  gmul3_3(83) <= to_unsigned(16#FC#, 8);
  gmul3_3(84) <= to_unsigned(16#FF#, 8);
  gmul3_3(85) <= to_unsigned(16#FA#, 8);
  gmul3_3(86) <= to_unsigned(16#F9#, 8);
  gmul3_3(87) <= to_unsigned(16#E8#, 8);
  gmul3_3(88) <= to_unsigned(16#EB#, 8);
  gmul3_3(89) <= to_unsigned(16#EE#, 8);
  gmul3_3(90) <= to_unsigned(16#ED#, 8);
  gmul3_3(91) <= to_unsigned(16#E4#, 8);
  gmul3_3(92) <= to_unsigned(16#E7#, 8);
  gmul3_3(93) <= to_unsigned(16#E2#, 8);
  gmul3_3(94) <= to_unsigned(16#E1#, 8);
  gmul3_3(95) <= to_unsigned(16#A0#, 8);
  gmul3_3(96) <= to_unsigned(16#A3#, 8);
  gmul3_3(97) <= to_unsigned(16#A6#, 8);
  gmul3_3(98) <= to_unsigned(16#A5#, 8);
  gmul3_3(99) <= to_unsigned(16#AC#, 8);
  gmul3_3(100) <= to_unsigned(16#AF#, 8);
  gmul3_3(101) <= to_unsigned(16#AA#, 8);
  gmul3_3(102) <= to_unsigned(16#A9#, 8);
  gmul3_3(103) <= to_unsigned(16#B8#, 8);
  gmul3_3(104) <= to_unsigned(16#BB#, 8);
  gmul3_3(105) <= to_unsigned(16#BE#, 8);
  gmul3_3(106) <= to_unsigned(16#BD#, 8);
  gmul3_3(107) <= to_unsigned(16#B4#, 8);
  gmul3_3(108) <= to_unsigned(16#B7#, 8);
  gmul3_3(109) <= to_unsigned(16#B2#, 8);
  gmul3_3(110) <= to_unsigned(16#B1#, 8);
  gmul3_3(111) <= to_unsigned(16#90#, 8);
  gmul3_3(112) <= to_unsigned(16#93#, 8);
  gmul3_3(113) <= to_unsigned(16#96#, 8);
  gmul3_3(114) <= to_unsigned(16#95#, 8);
  gmul3_3(115) <= to_unsigned(16#9C#, 8);
  gmul3_3(116) <= to_unsigned(16#9F#, 8);
  gmul3_3(117) <= to_unsigned(16#9A#, 8);
  gmul3_3(118) <= to_unsigned(16#99#, 8);
  gmul3_3(119) <= to_unsigned(16#88#, 8);
  gmul3_3(120) <= to_unsigned(16#8B#, 8);
  gmul3_3(121) <= to_unsigned(16#8E#, 8);
  gmul3_3(122) <= to_unsigned(16#8D#, 8);
  gmul3_3(123) <= to_unsigned(16#84#, 8);
  gmul3_3(124) <= to_unsigned(16#87#, 8);
  gmul3_3(125) <= to_unsigned(16#82#, 8);
  gmul3_3(126) <= to_unsigned(16#81#, 8);
  gmul3_3(127) <= to_unsigned(16#9B#, 8);
  gmul3_3(128) <= to_unsigned(16#98#, 8);
  gmul3_3(129) <= to_unsigned(16#9D#, 8);
  gmul3_3(130) <= to_unsigned(16#9E#, 8);
  gmul3_3(131) <= to_unsigned(16#97#, 8);
  gmul3_3(132) <= to_unsigned(16#94#, 8);
  gmul3_3(133) <= to_unsigned(16#91#, 8);
  gmul3_3(134) <= to_unsigned(16#92#, 8);
  gmul3_3(135) <= to_unsigned(16#83#, 8);
  gmul3_3(136) <= to_unsigned(16#80#, 8);
  gmul3_3(137) <= to_unsigned(16#85#, 8);
  gmul3_3(138) <= to_unsigned(16#86#, 8);
  gmul3_3(139) <= to_unsigned(16#8F#, 8);
  gmul3_3(140) <= to_unsigned(16#8C#, 8);
  gmul3_3(141) <= to_unsigned(16#89#, 8);
  gmul3_3(142) <= to_unsigned(16#8A#, 8);
  gmul3_3(143) <= to_unsigned(16#AB#, 8);
  gmul3_3(144) <= to_unsigned(16#A8#, 8);
  gmul3_3(145) <= to_unsigned(16#AD#, 8);
  gmul3_3(146) <= to_unsigned(16#AE#, 8);
  gmul3_3(147) <= to_unsigned(16#A7#, 8);
  gmul3_3(148) <= to_unsigned(16#A4#, 8);
  gmul3_3(149) <= to_unsigned(16#A1#, 8);
  gmul3_3(150) <= to_unsigned(16#A2#, 8);
  gmul3_3(151) <= to_unsigned(16#B3#, 8);
  gmul3_3(152) <= to_unsigned(16#B0#, 8);
  gmul3_3(153) <= to_unsigned(16#B5#, 8);
  gmul3_3(154) <= to_unsigned(16#B6#, 8);
  gmul3_3(155) <= to_unsigned(16#BF#, 8);
  gmul3_3(156) <= to_unsigned(16#BC#, 8);
  gmul3_3(157) <= to_unsigned(16#B9#, 8);
  gmul3_3(158) <= to_unsigned(16#BA#, 8);
  gmul3_3(159) <= to_unsigned(16#FB#, 8);
  gmul3_3(160) <= to_unsigned(16#F8#, 8);
  gmul3_3(161) <= to_unsigned(16#FD#, 8);
  gmul3_3(162) <= to_unsigned(16#FE#, 8);
  gmul3_3(163) <= to_unsigned(16#F7#, 8);
  gmul3_3(164) <= to_unsigned(16#F4#, 8);
  gmul3_3(165) <= to_unsigned(16#F1#, 8);
  gmul3_3(166) <= to_unsigned(16#F2#, 8);
  gmul3_3(167) <= to_unsigned(16#E3#, 8);
  gmul3_3(168) <= to_unsigned(16#E0#, 8);
  gmul3_3(169) <= to_unsigned(16#E5#, 8);
  gmul3_3(170) <= to_unsigned(16#E6#, 8);
  gmul3_3(171) <= to_unsigned(16#EF#, 8);
  gmul3_3(172) <= to_unsigned(16#EC#, 8);
  gmul3_3(173) <= to_unsigned(16#E9#, 8);
  gmul3_3(174) <= to_unsigned(16#EA#, 8);
  gmul3_3(175) <= to_unsigned(16#CB#, 8);
  gmul3_3(176) <= to_unsigned(16#C8#, 8);
  gmul3_3(177) <= to_unsigned(16#CD#, 8);
  gmul3_3(178) <= to_unsigned(16#CE#, 8);
  gmul3_3(179) <= to_unsigned(16#C7#, 8);
  gmul3_3(180) <= to_unsigned(16#C4#, 8);
  gmul3_3(181) <= to_unsigned(16#C1#, 8);
  gmul3_3(182) <= to_unsigned(16#C2#, 8);
  gmul3_3(183) <= to_unsigned(16#D3#, 8);
  gmul3_3(184) <= to_unsigned(16#D0#, 8);
  gmul3_3(185) <= to_unsigned(16#D5#, 8);
  gmul3_3(186) <= to_unsigned(16#D6#, 8);
  gmul3_3(187) <= to_unsigned(16#DF#, 8);
  gmul3_3(188) <= to_unsigned(16#DC#, 8);
  gmul3_3(189) <= to_unsigned(16#D9#, 8);
  gmul3_3(190) <= to_unsigned(16#DA#, 8);
  gmul3_3(191) <= to_unsigned(16#5B#, 8);
  gmul3_3(192) <= to_unsigned(16#58#, 8);
  gmul3_3(193) <= to_unsigned(16#5D#, 8);
  gmul3_3(194) <= to_unsigned(16#5E#, 8);
  gmul3_3(195) <= to_unsigned(16#57#, 8);
  gmul3_3(196) <= to_unsigned(16#54#, 8);
  gmul3_3(197) <= to_unsigned(16#51#, 8);
  gmul3_3(198) <= to_unsigned(16#52#, 8);
  gmul3_3(199) <= to_unsigned(16#43#, 8);
  gmul3_3(200) <= to_unsigned(16#40#, 8);
  gmul3_3(201) <= to_unsigned(16#45#, 8);
  gmul3_3(202) <= to_unsigned(16#46#, 8);
  gmul3_3(203) <= to_unsigned(16#4F#, 8);
  gmul3_3(204) <= to_unsigned(16#4C#, 8);
  gmul3_3(205) <= to_unsigned(16#49#, 8);
  gmul3_3(206) <= to_unsigned(16#4A#, 8);
  gmul3_3(207) <= to_unsigned(16#6B#, 8);
  gmul3_3(208) <= to_unsigned(16#68#, 8);
  gmul3_3(209) <= to_unsigned(16#6D#, 8);
  gmul3_3(210) <= to_unsigned(16#6E#, 8);
  gmul3_3(211) <= to_unsigned(16#67#, 8);
  gmul3_3(212) <= to_unsigned(16#64#, 8);
  gmul3_3(213) <= to_unsigned(16#61#, 8);
  gmul3_3(214) <= to_unsigned(16#62#, 8);
  gmul3_3(215) <= to_unsigned(16#73#, 8);
  gmul3_3(216) <= to_unsigned(16#70#, 8);
  gmul3_3(217) <= to_unsigned(16#75#, 8);
  gmul3_3(218) <= to_unsigned(16#76#, 8);
  gmul3_3(219) <= to_unsigned(16#7F#, 8);
  gmul3_3(220) <= to_unsigned(16#7C#, 8);
  gmul3_3(221) <= to_unsigned(16#79#, 8);
  gmul3_3(222) <= to_unsigned(16#7A#, 8);
  gmul3_3(223) <= to_unsigned(16#3B#, 8);
  gmul3_3(224) <= to_unsigned(16#38#, 8);
  gmul3_3(225) <= to_unsigned(16#3D#, 8);
  gmul3_3(226) <= to_unsigned(16#3E#, 8);
  gmul3_3(227) <= to_unsigned(16#37#, 8);
  gmul3_3(228) <= to_unsigned(16#34#, 8);
  gmul3_3(229) <= to_unsigned(16#31#, 8);
  gmul3_3(230) <= to_unsigned(16#32#, 8);
  gmul3_3(231) <= to_unsigned(16#23#, 8);
  gmul3_3(232) <= to_unsigned(16#20#, 8);
  gmul3_3(233) <= to_unsigned(16#25#, 8);
  gmul3_3(234) <= to_unsigned(16#26#, 8);
  gmul3_3(235) <= to_unsigned(16#2F#, 8);
  gmul3_3(236) <= to_unsigned(16#2C#, 8);
  gmul3_3(237) <= to_unsigned(16#29#, 8);
  gmul3_3(238) <= to_unsigned(16#2A#, 8);
  gmul3_3(239) <= to_unsigned(16#0B#, 8);
  gmul3_3(240) <= to_unsigned(16#08#, 8);
  gmul3_3(241) <= to_unsigned(16#0D#, 8);
  gmul3_3(242) <= to_unsigned(16#0E#, 8);
  gmul3_3(243) <= to_unsigned(16#07#, 8);
  gmul3_3(244) <= to_unsigned(16#04#, 8);
  gmul3_3(245) <= to_unsigned(16#01#, 8);
  gmul3_3(246) <= to_unsigned(16#02#, 8);
  gmul3_3(247) <= to_unsigned(16#13#, 8);
  gmul3_3(248) <= to_unsigned(16#10#, 8);
  gmul3_3(249) <= to_unsigned(16#15#, 8);
  gmul3_3(250) <= to_unsigned(16#16#, 8);
  gmul3_3(251) <= to_unsigned(16#1F#, 8);
  gmul3_3(252) <= to_unsigned(16#1C#, 8);
  gmul3_3(253) <= to_unsigned(16#19#, 8);
  gmul3_3(254) <= to_unsigned(16#1A#, 8);
  gmul3_3(255) <= to_unsigned(16#1A#, 8);

  gmul2_3(0) <= to_unsigned(16#02#, 8);
  gmul2_3(1) <= to_unsigned(16#04#, 8);
  gmul2_3(2) <= to_unsigned(16#06#, 8);
  gmul2_3(3) <= to_unsigned(16#08#, 8);
  gmul2_3(4) <= to_unsigned(16#0A#, 8);
  gmul2_3(5) <= to_unsigned(16#0C#, 8);
  gmul2_3(6) <= to_unsigned(16#0E#, 8);
  gmul2_3(7) <= to_unsigned(16#10#, 8);
  gmul2_3(8) <= to_unsigned(16#12#, 8);
  gmul2_3(9) <= to_unsigned(16#14#, 8);
  gmul2_3(10) <= to_unsigned(16#16#, 8);
  gmul2_3(11) <= to_unsigned(16#18#, 8);
  gmul2_3(12) <= to_unsigned(16#1A#, 8);
  gmul2_3(13) <= to_unsigned(16#1C#, 8);
  gmul2_3(14) <= to_unsigned(16#1E#, 8);
  gmul2_3(15) <= to_unsigned(16#20#, 8);
  gmul2_3(16) <= to_unsigned(16#22#, 8);
  gmul2_3(17) <= to_unsigned(16#24#, 8);
  gmul2_3(18) <= to_unsigned(16#26#, 8);
  gmul2_3(19) <= to_unsigned(16#28#, 8);
  gmul2_3(20) <= to_unsigned(16#2A#, 8);
  gmul2_3(21) <= to_unsigned(16#2C#, 8);
  gmul2_3(22) <= to_unsigned(16#2E#, 8);
  gmul2_3(23) <= to_unsigned(16#30#, 8);
  gmul2_3(24) <= to_unsigned(16#32#, 8);
  gmul2_3(25) <= to_unsigned(16#34#, 8);
  gmul2_3(26) <= to_unsigned(16#36#, 8);
  gmul2_3(27) <= to_unsigned(16#38#, 8);
  gmul2_3(28) <= to_unsigned(16#3A#, 8);
  gmul2_3(29) <= to_unsigned(16#3C#, 8);
  gmul2_3(30) <= to_unsigned(16#3E#, 8);
  gmul2_3(31) <= to_unsigned(16#40#, 8);
  gmul2_3(32) <= to_unsigned(16#42#, 8);
  gmul2_3(33) <= to_unsigned(16#44#, 8);
  gmul2_3(34) <= to_unsigned(16#46#, 8);
  gmul2_3(35) <= to_unsigned(16#48#, 8);
  gmul2_3(36) <= to_unsigned(16#4A#, 8);
  gmul2_3(37) <= to_unsigned(16#4C#, 8);
  gmul2_3(38) <= to_unsigned(16#4E#, 8);
  gmul2_3(39) <= to_unsigned(16#50#, 8);
  gmul2_3(40) <= to_unsigned(16#52#, 8);
  gmul2_3(41) <= to_unsigned(16#54#, 8);
  gmul2_3(42) <= to_unsigned(16#56#, 8);
  gmul2_3(43) <= to_unsigned(16#58#, 8);
  gmul2_3(44) <= to_unsigned(16#5A#, 8);
  gmul2_3(45) <= to_unsigned(16#5C#, 8);
  gmul2_3(46) <= to_unsigned(16#5E#, 8);
  gmul2_3(47) <= to_unsigned(16#60#, 8);
  gmul2_3(48) <= to_unsigned(16#62#, 8);
  gmul2_3(49) <= to_unsigned(16#64#, 8);
  gmul2_3(50) <= to_unsigned(16#66#, 8);
  gmul2_3(51) <= to_unsigned(16#68#, 8);
  gmul2_3(52) <= to_unsigned(16#6A#, 8);
  gmul2_3(53) <= to_unsigned(16#6C#, 8);
  gmul2_3(54) <= to_unsigned(16#6E#, 8);
  gmul2_3(55) <= to_unsigned(16#70#, 8);
  gmul2_3(56) <= to_unsigned(16#72#, 8);
  gmul2_3(57) <= to_unsigned(16#74#, 8);
  gmul2_3(58) <= to_unsigned(16#76#, 8);
  gmul2_3(59) <= to_unsigned(16#78#, 8);
  gmul2_3(60) <= to_unsigned(16#7A#, 8);
  gmul2_3(61) <= to_unsigned(16#7C#, 8);
  gmul2_3(62) <= to_unsigned(16#7E#, 8);
  gmul2_3(63) <= to_unsigned(16#80#, 8);
  gmul2_3(64) <= to_unsigned(16#82#, 8);
  gmul2_3(65) <= to_unsigned(16#84#, 8);
  gmul2_3(66) <= to_unsigned(16#86#, 8);
  gmul2_3(67) <= to_unsigned(16#88#, 8);
  gmul2_3(68) <= to_unsigned(16#8A#, 8);
  gmul2_3(69) <= to_unsigned(16#8C#, 8);
  gmul2_3(70) <= to_unsigned(16#8E#, 8);
  gmul2_3(71) <= to_unsigned(16#90#, 8);
  gmul2_3(72) <= to_unsigned(16#92#, 8);
  gmul2_3(73) <= to_unsigned(16#94#, 8);
  gmul2_3(74) <= to_unsigned(16#96#, 8);
  gmul2_3(75) <= to_unsigned(16#98#, 8);
  gmul2_3(76) <= to_unsigned(16#9A#, 8);
  gmul2_3(77) <= to_unsigned(16#9C#, 8);
  gmul2_3(78) <= to_unsigned(16#9E#, 8);
  gmul2_3(79) <= to_unsigned(16#A0#, 8);
  gmul2_3(80) <= to_unsigned(16#A2#, 8);
  gmul2_3(81) <= to_unsigned(16#A4#, 8);
  gmul2_3(82) <= to_unsigned(16#A6#, 8);
  gmul2_3(83) <= to_unsigned(16#A8#, 8);
  gmul2_3(84) <= to_unsigned(16#AA#, 8);
  gmul2_3(85) <= to_unsigned(16#AC#, 8);
  gmul2_3(86) <= to_unsigned(16#AE#, 8);
  gmul2_3(87) <= to_unsigned(16#B0#, 8);
  gmul2_3(88) <= to_unsigned(16#B2#, 8);
  gmul2_3(89) <= to_unsigned(16#B4#, 8);
  gmul2_3(90) <= to_unsigned(16#B6#, 8);
  gmul2_3(91) <= to_unsigned(16#B8#, 8);
  gmul2_3(92) <= to_unsigned(16#BA#, 8);
  gmul2_3(93) <= to_unsigned(16#BC#, 8);
  gmul2_3(94) <= to_unsigned(16#BE#, 8);
  gmul2_3(95) <= to_unsigned(16#C0#, 8);
  gmul2_3(96) <= to_unsigned(16#C2#, 8);
  gmul2_3(97) <= to_unsigned(16#C4#, 8);
  gmul2_3(98) <= to_unsigned(16#C6#, 8);
  gmul2_3(99) <= to_unsigned(16#C8#, 8);
  gmul2_3(100) <= to_unsigned(16#CA#, 8);
  gmul2_3(101) <= to_unsigned(16#CC#, 8);
  gmul2_3(102) <= to_unsigned(16#CE#, 8);
  gmul2_3(103) <= to_unsigned(16#D0#, 8);
  gmul2_3(104) <= to_unsigned(16#D2#, 8);
  gmul2_3(105) <= to_unsigned(16#D4#, 8);
  gmul2_3(106) <= to_unsigned(16#D6#, 8);
  gmul2_3(107) <= to_unsigned(16#D8#, 8);
  gmul2_3(108) <= to_unsigned(16#DA#, 8);
  gmul2_3(109) <= to_unsigned(16#DC#, 8);
  gmul2_3(110) <= to_unsigned(16#DE#, 8);
  gmul2_3(111) <= to_unsigned(16#E0#, 8);
  gmul2_3(112) <= to_unsigned(16#E2#, 8);
  gmul2_3(113) <= to_unsigned(16#E4#, 8);
  gmul2_3(114) <= to_unsigned(16#E6#, 8);
  gmul2_3(115) <= to_unsigned(16#E8#, 8);
  gmul2_3(116) <= to_unsigned(16#EA#, 8);
  gmul2_3(117) <= to_unsigned(16#EC#, 8);
  gmul2_3(118) <= to_unsigned(16#EE#, 8);
  gmul2_3(119) <= to_unsigned(16#F0#, 8);
  gmul2_3(120) <= to_unsigned(16#F2#, 8);
  gmul2_3(121) <= to_unsigned(16#F4#, 8);
  gmul2_3(122) <= to_unsigned(16#F6#, 8);
  gmul2_3(123) <= to_unsigned(16#F8#, 8);
  gmul2_3(124) <= to_unsigned(16#FA#, 8);
  gmul2_3(125) <= to_unsigned(16#FC#, 8);
  gmul2_3(126) <= to_unsigned(16#FE#, 8);
  gmul2_3(127) <= to_unsigned(16#1B#, 8);
  gmul2_3(128) <= to_unsigned(16#19#, 8);
  gmul2_3(129) <= to_unsigned(16#1F#, 8);
  gmul2_3(130) <= to_unsigned(16#1D#, 8);
  gmul2_3(131) <= to_unsigned(16#13#, 8);
  gmul2_3(132) <= to_unsigned(16#11#, 8);
  gmul2_3(133) <= to_unsigned(16#17#, 8);
  gmul2_3(134) <= to_unsigned(16#15#, 8);
  gmul2_3(135) <= to_unsigned(16#0B#, 8);
  gmul2_3(136) <= to_unsigned(16#09#, 8);
  gmul2_3(137) <= to_unsigned(16#0F#, 8);
  gmul2_3(138) <= to_unsigned(16#0D#, 8);
  gmul2_3(139) <= to_unsigned(16#03#, 8);
  gmul2_3(140) <= to_unsigned(16#01#, 8);
  gmul2_3(141) <= to_unsigned(16#07#, 8);
  gmul2_3(142) <= to_unsigned(16#05#, 8);
  gmul2_3(143) <= to_unsigned(16#3B#, 8);
  gmul2_3(144) <= to_unsigned(16#39#, 8);
  gmul2_3(145) <= to_unsigned(16#3F#, 8);
  gmul2_3(146) <= to_unsigned(16#3D#, 8);
  gmul2_3(147) <= to_unsigned(16#33#, 8);
  gmul2_3(148) <= to_unsigned(16#31#, 8);
  gmul2_3(149) <= to_unsigned(16#37#, 8);
  gmul2_3(150) <= to_unsigned(16#35#, 8);
  gmul2_3(151) <= to_unsigned(16#2B#, 8);
  gmul2_3(152) <= to_unsigned(16#29#, 8);
  gmul2_3(153) <= to_unsigned(16#2F#, 8);
  gmul2_3(154) <= to_unsigned(16#2D#, 8);
  gmul2_3(155) <= to_unsigned(16#23#, 8);
  gmul2_3(156) <= to_unsigned(16#21#, 8);
  gmul2_3(157) <= to_unsigned(16#27#, 8);
  gmul2_3(158) <= to_unsigned(16#25#, 8);
  gmul2_3(159) <= to_unsigned(16#5B#, 8);
  gmul2_3(160) <= to_unsigned(16#59#, 8);
  gmul2_3(161) <= to_unsigned(16#5F#, 8);
  gmul2_3(162) <= to_unsigned(16#5D#, 8);
  gmul2_3(163) <= to_unsigned(16#53#, 8);
  gmul2_3(164) <= to_unsigned(16#51#, 8);
  gmul2_3(165) <= to_unsigned(16#57#, 8);
  gmul2_3(166) <= to_unsigned(16#55#, 8);
  gmul2_3(167) <= to_unsigned(16#4B#, 8);
  gmul2_3(168) <= to_unsigned(16#49#, 8);
  gmul2_3(169) <= to_unsigned(16#4F#, 8);
  gmul2_3(170) <= to_unsigned(16#4D#, 8);
  gmul2_3(171) <= to_unsigned(16#43#, 8);
  gmul2_3(172) <= to_unsigned(16#41#, 8);
  gmul2_3(173) <= to_unsigned(16#47#, 8);
  gmul2_3(174) <= to_unsigned(16#45#, 8);
  gmul2_3(175) <= to_unsigned(16#7B#, 8);
  gmul2_3(176) <= to_unsigned(16#79#, 8);
  gmul2_3(177) <= to_unsigned(16#7F#, 8);
  gmul2_3(178) <= to_unsigned(16#7D#, 8);
  gmul2_3(179) <= to_unsigned(16#73#, 8);
  gmul2_3(180) <= to_unsigned(16#71#, 8);
  gmul2_3(181) <= to_unsigned(16#77#, 8);
  gmul2_3(182) <= to_unsigned(16#75#, 8);
  gmul2_3(183) <= to_unsigned(16#6B#, 8);
  gmul2_3(184) <= to_unsigned(16#69#, 8);
  gmul2_3(185) <= to_unsigned(16#6F#, 8);
  gmul2_3(186) <= to_unsigned(16#6D#, 8);
  gmul2_3(187) <= to_unsigned(16#63#, 8);
  gmul2_3(188) <= to_unsigned(16#61#, 8);
  gmul2_3(189) <= to_unsigned(16#67#, 8);
  gmul2_3(190) <= to_unsigned(16#65#, 8);
  gmul2_3(191) <= to_unsigned(16#9B#, 8);
  gmul2_3(192) <= to_unsigned(16#99#, 8);
  gmul2_3(193) <= to_unsigned(16#9F#, 8);
  gmul2_3(194) <= to_unsigned(16#9D#, 8);
  gmul2_3(195) <= to_unsigned(16#93#, 8);
  gmul2_3(196) <= to_unsigned(16#91#, 8);
  gmul2_3(197) <= to_unsigned(16#97#, 8);
  gmul2_3(198) <= to_unsigned(16#95#, 8);
  gmul2_3(199) <= to_unsigned(16#8B#, 8);
  gmul2_3(200) <= to_unsigned(16#89#, 8);
  gmul2_3(201) <= to_unsigned(16#8F#, 8);
  gmul2_3(202) <= to_unsigned(16#8D#, 8);
  gmul2_3(203) <= to_unsigned(16#83#, 8);
  gmul2_3(204) <= to_unsigned(16#81#, 8);
  gmul2_3(205) <= to_unsigned(16#87#, 8);
  gmul2_3(206) <= to_unsigned(16#85#, 8);
  gmul2_3(207) <= to_unsigned(16#BB#, 8);
  gmul2_3(208) <= to_unsigned(16#B9#, 8);
  gmul2_3(209) <= to_unsigned(16#BF#, 8);
  gmul2_3(210) <= to_unsigned(16#BD#, 8);
  gmul2_3(211) <= to_unsigned(16#B3#, 8);
  gmul2_3(212) <= to_unsigned(16#B1#, 8);
  gmul2_3(213) <= to_unsigned(16#B7#, 8);
  gmul2_3(214) <= to_unsigned(16#B5#, 8);
  gmul2_3(215) <= to_unsigned(16#AB#, 8);
  gmul2_3(216) <= to_unsigned(16#A9#, 8);
  gmul2_3(217) <= to_unsigned(16#AF#, 8);
  gmul2_3(218) <= to_unsigned(16#AD#, 8);
  gmul2_3(219) <= to_unsigned(16#A3#, 8);
  gmul2_3(220) <= to_unsigned(16#A1#, 8);
  gmul2_3(221) <= to_unsigned(16#A7#, 8);
  gmul2_3(222) <= to_unsigned(16#A5#, 8);
  gmul2_3(223) <= to_unsigned(16#DB#, 8);
  gmul2_3(224) <= to_unsigned(16#D9#, 8);
  gmul2_3(225) <= to_unsigned(16#DF#, 8);
  gmul2_3(226) <= to_unsigned(16#DD#, 8);
  gmul2_3(227) <= to_unsigned(16#D3#, 8);
  gmul2_3(228) <= to_unsigned(16#D1#, 8);
  gmul2_3(229) <= to_unsigned(16#D7#, 8);
  gmul2_3(230) <= to_unsigned(16#D5#, 8);
  gmul2_3(231) <= to_unsigned(16#CB#, 8);
  gmul2_3(232) <= to_unsigned(16#C9#, 8);
  gmul2_3(233) <= to_unsigned(16#CF#, 8);
  gmul2_3(234) <= to_unsigned(16#CD#, 8);
  gmul2_3(235) <= to_unsigned(16#C3#, 8);
  gmul2_3(236) <= to_unsigned(16#C1#, 8);
  gmul2_3(237) <= to_unsigned(16#C7#, 8);
  gmul2_3(238) <= to_unsigned(16#C5#, 8);
  gmul2_3(239) <= to_unsigned(16#FB#, 8);
  gmul2_3(240) <= to_unsigned(16#F9#, 8);
  gmul2_3(241) <= to_unsigned(16#FF#, 8);
  gmul2_3(242) <= to_unsigned(16#FD#, 8);
  gmul2_3(243) <= to_unsigned(16#F3#, 8);
  gmul2_3(244) <= to_unsigned(16#F1#, 8);
  gmul2_3(245) <= to_unsigned(16#F7#, 8);
  gmul2_3(246) <= to_unsigned(16#F5#, 8);
  gmul2_3(247) <= to_unsigned(16#EB#, 8);
  gmul2_3(248) <= to_unsigned(16#E9#, 8);
  gmul2_3(249) <= to_unsigned(16#EF#, 8);
  gmul2_3(250) <= to_unsigned(16#ED#, 8);
  gmul2_3(251) <= to_unsigned(16#E3#, 8);
  gmul2_3(252) <= to_unsigned(16#E1#, 8);
  gmul2_3(253) <= to_unsigned(16#E7#, 8);
  gmul2_3(254) <= to_unsigned(16#E5#, 8);
  gmul2_3(255) <= to_unsigned(16#E5#, 8);

  gmul2_4(0) <= to_unsigned(16#02#, 8);
  gmul2_4(1) <= to_unsigned(16#04#, 8);
  gmul2_4(2) <= to_unsigned(16#06#, 8);
  gmul2_4(3) <= to_unsigned(16#08#, 8);
  gmul2_4(4) <= to_unsigned(16#0A#, 8);
  gmul2_4(5) <= to_unsigned(16#0C#, 8);
  gmul2_4(6) <= to_unsigned(16#0E#, 8);
  gmul2_4(7) <= to_unsigned(16#10#, 8);
  gmul2_4(8) <= to_unsigned(16#12#, 8);
  gmul2_4(9) <= to_unsigned(16#14#, 8);
  gmul2_4(10) <= to_unsigned(16#16#, 8);
  gmul2_4(11) <= to_unsigned(16#18#, 8);
  gmul2_4(12) <= to_unsigned(16#1A#, 8);
  gmul2_4(13) <= to_unsigned(16#1C#, 8);
  gmul2_4(14) <= to_unsigned(16#1E#, 8);
  gmul2_4(15) <= to_unsigned(16#20#, 8);
  gmul2_4(16) <= to_unsigned(16#22#, 8);
  gmul2_4(17) <= to_unsigned(16#24#, 8);
  gmul2_4(18) <= to_unsigned(16#26#, 8);
  gmul2_4(19) <= to_unsigned(16#28#, 8);
  gmul2_4(20) <= to_unsigned(16#2A#, 8);
  gmul2_4(21) <= to_unsigned(16#2C#, 8);
  gmul2_4(22) <= to_unsigned(16#2E#, 8);
  gmul2_4(23) <= to_unsigned(16#30#, 8);
  gmul2_4(24) <= to_unsigned(16#32#, 8);
  gmul2_4(25) <= to_unsigned(16#34#, 8);
  gmul2_4(26) <= to_unsigned(16#36#, 8);
  gmul2_4(27) <= to_unsigned(16#38#, 8);
  gmul2_4(28) <= to_unsigned(16#3A#, 8);
  gmul2_4(29) <= to_unsigned(16#3C#, 8);
  gmul2_4(30) <= to_unsigned(16#3E#, 8);
  gmul2_4(31) <= to_unsigned(16#40#, 8);
  gmul2_4(32) <= to_unsigned(16#42#, 8);
  gmul2_4(33) <= to_unsigned(16#44#, 8);
  gmul2_4(34) <= to_unsigned(16#46#, 8);
  gmul2_4(35) <= to_unsigned(16#48#, 8);
  gmul2_4(36) <= to_unsigned(16#4A#, 8);
  gmul2_4(37) <= to_unsigned(16#4C#, 8);
  gmul2_4(38) <= to_unsigned(16#4E#, 8);
  gmul2_4(39) <= to_unsigned(16#50#, 8);
  gmul2_4(40) <= to_unsigned(16#52#, 8);
  gmul2_4(41) <= to_unsigned(16#54#, 8);
  gmul2_4(42) <= to_unsigned(16#56#, 8);
  gmul2_4(43) <= to_unsigned(16#58#, 8);
  gmul2_4(44) <= to_unsigned(16#5A#, 8);
  gmul2_4(45) <= to_unsigned(16#5C#, 8);
  gmul2_4(46) <= to_unsigned(16#5E#, 8);
  gmul2_4(47) <= to_unsigned(16#60#, 8);
  gmul2_4(48) <= to_unsigned(16#62#, 8);
  gmul2_4(49) <= to_unsigned(16#64#, 8);
  gmul2_4(50) <= to_unsigned(16#66#, 8);
  gmul2_4(51) <= to_unsigned(16#68#, 8);
  gmul2_4(52) <= to_unsigned(16#6A#, 8);
  gmul2_4(53) <= to_unsigned(16#6C#, 8);
  gmul2_4(54) <= to_unsigned(16#6E#, 8);
  gmul2_4(55) <= to_unsigned(16#70#, 8);
  gmul2_4(56) <= to_unsigned(16#72#, 8);
  gmul2_4(57) <= to_unsigned(16#74#, 8);
  gmul2_4(58) <= to_unsigned(16#76#, 8);
  gmul2_4(59) <= to_unsigned(16#78#, 8);
  gmul2_4(60) <= to_unsigned(16#7A#, 8);
  gmul2_4(61) <= to_unsigned(16#7C#, 8);
  gmul2_4(62) <= to_unsigned(16#7E#, 8);
  gmul2_4(63) <= to_unsigned(16#80#, 8);
  gmul2_4(64) <= to_unsigned(16#82#, 8);
  gmul2_4(65) <= to_unsigned(16#84#, 8);
  gmul2_4(66) <= to_unsigned(16#86#, 8);
  gmul2_4(67) <= to_unsigned(16#88#, 8);
  gmul2_4(68) <= to_unsigned(16#8A#, 8);
  gmul2_4(69) <= to_unsigned(16#8C#, 8);
  gmul2_4(70) <= to_unsigned(16#8E#, 8);
  gmul2_4(71) <= to_unsigned(16#90#, 8);
  gmul2_4(72) <= to_unsigned(16#92#, 8);
  gmul2_4(73) <= to_unsigned(16#94#, 8);
  gmul2_4(74) <= to_unsigned(16#96#, 8);
  gmul2_4(75) <= to_unsigned(16#98#, 8);
  gmul2_4(76) <= to_unsigned(16#9A#, 8);
  gmul2_4(77) <= to_unsigned(16#9C#, 8);
  gmul2_4(78) <= to_unsigned(16#9E#, 8);
  gmul2_4(79) <= to_unsigned(16#A0#, 8);
  gmul2_4(80) <= to_unsigned(16#A2#, 8);
  gmul2_4(81) <= to_unsigned(16#A4#, 8);
  gmul2_4(82) <= to_unsigned(16#A6#, 8);
  gmul2_4(83) <= to_unsigned(16#A8#, 8);
  gmul2_4(84) <= to_unsigned(16#AA#, 8);
  gmul2_4(85) <= to_unsigned(16#AC#, 8);
  gmul2_4(86) <= to_unsigned(16#AE#, 8);
  gmul2_4(87) <= to_unsigned(16#B0#, 8);
  gmul2_4(88) <= to_unsigned(16#B2#, 8);
  gmul2_4(89) <= to_unsigned(16#B4#, 8);
  gmul2_4(90) <= to_unsigned(16#B6#, 8);
  gmul2_4(91) <= to_unsigned(16#B8#, 8);
  gmul2_4(92) <= to_unsigned(16#BA#, 8);
  gmul2_4(93) <= to_unsigned(16#BC#, 8);
  gmul2_4(94) <= to_unsigned(16#BE#, 8);
  gmul2_4(95) <= to_unsigned(16#C0#, 8);
  gmul2_4(96) <= to_unsigned(16#C2#, 8);
  gmul2_4(97) <= to_unsigned(16#C4#, 8);
  gmul2_4(98) <= to_unsigned(16#C6#, 8);
  gmul2_4(99) <= to_unsigned(16#C8#, 8);
  gmul2_4(100) <= to_unsigned(16#CA#, 8);
  gmul2_4(101) <= to_unsigned(16#CC#, 8);
  gmul2_4(102) <= to_unsigned(16#CE#, 8);
  gmul2_4(103) <= to_unsigned(16#D0#, 8);
  gmul2_4(104) <= to_unsigned(16#D2#, 8);
  gmul2_4(105) <= to_unsigned(16#D4#, 8);
  gmul2_4(106) <= to_unsigned(16#D6#, 8);
  gmul2_4(107) <= to_unsigned(16#D8#, 8);
  gmul2_4(108) <= to_unsigned(16#DA#, 8);
  gmul2_4(109) <= to_unsigned(16#DC#, 8);
  gmul2_4(110) <= to_unsigned(16#DE#, 8);
  gmul2_4(111) <= to_unsigned(16#E0#, 8);
  gmul2_4(112) <= to_unsigned(16#E2#, 8);
  gmul2_4(113) <= to_unsigned(16#E4#, 8);
  gmul2_4(114) <= to_unsigned(16#E6#, 8);
  gmul2_4(115) <= to_unsigned(16#E8#, 8);
  gmul2_4(116) <= to_unsigned(16#EA#, 8);
  gmul2_4(117) <= to_unsigned(16#EC#, 8);
  gmul2_4(118) <= to_unsigned(16#EE#, 8);
  gmul2_4(119) <= to_unsigned(16#F0#, 8);
  gmul2_4(120) <= to_unsigned(16#F2#, 8);
  gmul2_4(121) <= to_unsigned(16#F4#, 8);
  gmul2_4(122) <= to_unsigned(16#F6#, 8);
  gmul2_4(123) <= to_unsigned(16#F8#, 8);
  gmul2_4(124) <= to_unsigned(16#FA#, 8);
  gmul2_4(125) <= to_unsigned(16#FC#, 8);
  gmul2_4(126) <= to_unsigned(16#FE#, 8);
  gmul2_4(127) <= to_unsigned(16#1B#, 8);
  gmul2_4(128) <= to_unsigned(16#19#, 8);
  gmul2_4(129) <= to_unsigned(16#1F#, 8);
  gmul2_4(130) <= to_unsigned(16#1D#, 8);
  gmul2_4(131) <= to_unsigned(16#13#, 8);
  gmul2_4(132) <= to_unsigned(16#11#, 8);
  gmul2_4(133) <= to_unsigned(16#17#, 8);
  gmul2_4(134) <= to_unsigned(16#15#, 8);
  gmul2_4(135) <= to_unsigned(16#0B#, 8);
  gmul2_4(136) <= to_unsigned(16#09#, 8);
  gmul2_4(137) <= to_unsigned(16#0F#, 8);
  gmul2_4(138) <= to_unsigned(16#0D#, 8);
  gmul2_4(139) <= to_unsigned(16#03#, 8);
  gmul2_4(140) <= to_unsigned(16#01#, 8);
  gmul2_4(141) <= to_unsigned(16#07#, 8);
  gmul2_4(142) <= to_unsigned(16#05#, 8);
  gmul2_4(143) <= to_unsigned(16#3B#, 8);
  gmul2_4(144) <= to_unsigned(16#39#, 8);
  gmul2_4(145) <= to_unsigned(16#3F#, 8);
  gmul2_4(146) <= to_unsigned(16#3D#, 8);
  gmul2_4(147) <= to_unsigned(16#33#, 8);
  gmul2_4(148) <= to_unsigned(16#31#, 8);
  gmul2_4(149) <= to_unsigned(16#37#, 8);
  gmul2_4(150) <= to_unsigned(16#35#, 8);
  gmul2_4(151) <= to_unsigned(16#2B#, 8);
  gmul2_4(152) <= to_unsigned(16#29#, 8);
  gmul2_4(153) <= to_unsigned(16#2F#, 8);
  gmul2_4(154) <= to_unsigned(16#2D#, 8);
  gmul2_4(155) <= to_unsigned(16#23#, 8);
  gmul2_4(156) <= to_unsigned(16#21#, 8);
  gmul2_4(157) <= to_unsigned(16#27#, 8);
  gmul2_4(158) <= to_unsigned(16#25#, 8);
  gmul2_4(159) <= to_unsigned(16#5B#, 8);
  gmul2_4(160) <= to_unsigned(16#59#, 8);
  gmul2_4(161) <= to_unsigned(16#5F#, 8);
  gmul2_4(162) <= to_unsigned(16#5D#, 8);
  gmul2_4(163) <= to_unsigned(16#53#, 8);
  gmul2_4(164) <= to_unsigned(16#51#, 8);
  gmul2_4(165) <= to_unsigned(16#57#, 8);
  gmul2_4(166) <= to_unsigned(16#55#, 8);
  gmul2_4(167) <= to_unsigned(16#4B#, 8);
  gmul2_4(168) <= to_unsigned(16#49#, 8);
  gmul2_4(169) <= to_unsigned(16#4F#, 8);
  gmul2_4(170) <= to_unsigned(16#4D#, 8);
  gmul2_4(171) <= to_unsigned(16#43#, 8);
  gmul2_4(172) <= to_unsigned(16#41#, 8);
  gmul2_4(173) <= to_unsigned(16#47#, 8);
  gmul2_4(174) <= to_unsigned(16#45#, 8);
  gmul2_4(175) <= to_unsigned(16#7B#, 8);
  gmul2_4(176) <= to_unsigned(16#79#, 8);
  gmul2_4(177) <= to_unsigned(16#7F#, 8);
  gmul2_4(178) <= to_unsigned(16#7D#, 8);
  gmul2_4(179) <= to_unsigned(16#73#, 8);
  gmul2_4(180) <= to_unsigned(16#71#, 8);
  gmul2_4(181) <= to_unsigned(16#77#, 8);
  gmul2_4(182) <= to_unsigned(16#75#, 8);
  gmul2_4(183) <= to_unsigned(16#6B#, 8);
  gmul2_4(184) <= to_unsigned(16#69#, 8);
  gmul2_4(185) <= to_unsigned(16#6F#, 8);
  gmul2_4(186) <= to_unsigned(16#6D#, 8);
  gmul2_4(187) <= to_unsigned(16#63#, 8);
  gmul2_4(188) <= to_unsigned(16#61#, 8);
  gmul2_4(189) <= to_unsigned(16#67#, 8);
  gmul2_4(190) <= to_unsigned(16#65#, 8);
  gmul2_4(191) <= to_unsigned(16#9B#, 8);
  gmul2_4(192) <= to_unsigned(16#99#, 8);
  gmul2_4(193) <= to_unsigned(16#9F#, 8);
  gmul2_4(194) <= to_unsigned(16#9D#, 8);
  gmul2_4(195) <= to_unsigned(16#93#, 8);
  gmul2_4(196) <= to_unsigned(16#91#, 8);
  gmul2_4(197) <= to_unsigned(16#97#, 8);
  gmul2_4(198) <= to_unsigned(16#95#, 8);
  gmul2_4(199) <= to_unsigned(16#8B#, 8);
  gmul2_4(200) <= to_unsigned(16#89#, 8);
  gmul2_4(201) <= to_unsigned(16#8F#, 8);
  gmul2_4(202) <= to_unsigned(16#8D#, 8);
  gmul2_4(203) <= to_unsigned(16#83#, 8);
  gmul2_4(204) <= to_unsigned(16#81#, 8);
  gmul2_4(205) <= to_unsigned(16#87#, 8);
  gmul2_4(206) <= to_unsigned(16#85#, 8);
  gmul2_4(207) <= to_unsigned(16#BB#, 8);
  gmul2_4(208) <= to_unsigned(16#B9#, 8);
  gmul2_4(209) <= to_unsigned(16#BF#, 8);
  gmul2_4(210) <= to_unsigned(16#BD#, 8);
  gmul2_4(211) <= to_unsigned(16#B3#, 8);
  gmul2_4(212) <= to_unsigned(16#B1#, 8);
  gmul2_4(213) <= to_unsigned(16#B7#, 8);
  gmul2_4(214) <= to_unsigned(16#B5#, 8);
  gmul2_4(215) <= to_unsigned(16#AB#, 8);
  gmul2_4(216) <= to_unsigned(16#A9#, 8);
  gmul2_4(217) <= to_unsigned(16#AF#, 8);
  gmul2_4(218) <= to_unsigned(16#AD#, 8);
  gmul2_4(219) <= to_unsigned(16#A3#, 8);
  gmul2_4(220) <= to_unsigned(16#A1#, 8);
  gmul2_4(221) <= to_unsigned(16#A7#, 8);
  gmul2_4(222) <= to_unsigned(16#A5#, 8);
  gmul2_4(223) <= to_unsigned(16#DB#, 8);
  gmul2_4(224) <= to_unsigned(16#D9#, 8);
  gmul2_4(225) <= to_unsigned(16#DF#, 8);
  gmul2_4(226) <= to_unsigned(16#DD#, 8);
  gmul2_4(227) <= to_unsigned(16#D3#, 8);
  gmul2_4(228) <= to_unsigned(16#D1#, 8);
  gmul2_4(229) <= to_unsigned(16#D7#, 8);
  gmul2_4(230) <= to_unsigned(16#D5#, 8);
  gmul2_4(231) <= to_unsigned(16#CB#, 8);
  gmul2_4(232) <= to_unsigned(16#C9#, 8);
  gmul2_4(233) <= to_unsigned(16#CF#, 8);
  gmul2_4(234) <= to_unsigned(16#CD#, 8);
  gmul2_4(235) <= to_unsigned(16#C3#, 8);
  gmul2_4(236) <= to_unsigned(16#C1#, 8);
  gmul2_4(237) <= to_unsigned(16#C7#, 8);
  gmul2_4(238) <= to_unsigned(16#C5#, 8);
  gmul2_4(239) <= to_unsigned(16#FB#, 8);
  gmul2_4(240) <= to_unsigned(16#F9#, 8);
  gmul2_4(241) <= to_unsigned(16#FF#, 8);
  gmul2_4(242) <= to_unsigned(16#FD#, 8);
  gmul2_4(243) <= to_unsigned(16#F3#, 8);
  gmul2_4(244) <= to_unsigned(16#F1#, 8);
  gmul2_4(245) <= to_unsigned(16#F7#, 8);
  gmul2_4(246) <= to_unsigned(16#F5#, 8);
  gmul2_4(247) <= to_unsigned(16#EB#, 8);
  gmul2_4(248) <= to_unsigned(16#E9#, 8);
  gmul2_4(249) <= to_unsigned(16#EF#, 8);
  gmul2_4(250) <= to_unsigned(16#ED#, 8);
  gmul2_4(251) <= to_unsigned(16#E3#, 8);
  gmul2_4(252) <= to_unsigned(16#E1#, 8);
  gmul2_4(253) <= to_unsigned(16#E7#, 8);
  gmul2_4(254) <= to_unsigned(16#E5#, 8);
  gmul2_4(255) <= to_unsigned(16#E5#, 8);

  gmul3_4(0) <= to_unsigned(16#03#, 8);
  gmul3_4(1) <= to_unsigned(16#06#, 8);
  gmul3_4(2) <= to_unsigned(16#05#, 8);
  gmul3_4(3) <= to_unsigned(16#0C#, 8);
  gmul3_4(4) <= to_unsigned(16#0F#, 8);
  gmul3_4(5) <= to_unsigned(16#0A#, 8);
  gmul3_4(6) <= to_unsigned(16#09#, 8);
  gmul3_4(7) <= to_unsigned(16#18#, 8);
  gmul3_4(8) <= to_unsigned(16#1B#, 8);
  gmul3_4(9) <= to_unsigned(16#1E#, 8);
  gmul3_4(10) <= to_unsigned(16#1D#, 8);
  gmul3_4(11) <= to_unsigned(16#14#, 8);
  gmul3_4(12) <= to_unsigned(16#17#, 8);
  gmul3_4(13) <= to_unsigned(16#12#, 8);
  gmul3_4(14) <= to_unsigned(16#11#, 8);
  gmul3_4(15) <= to_unsigned(16#30#, 8);
  gmul3_4(16) <= to_unsigned(16#33#, 8);
  gmul3_4(17) <= to_unsigned(16#36#, 8);
  gmul3_4(18) <= to_unsigned(16#35#, 8);
  gmul3_4(19) <= to_unsigned(16#3C#, 8);
  gmul3_4(20) <= to_unsigned(16#3F#, 8);
  gmul3_4(21) <= to_unsigned(16#3A#, 8);
  gmul3_4(22) <= to_unsigned(16#39#, 8);
  gmul3_4(23) <= to_unsigned(16#28#, 8);
  gmul3_4(24) <= to_unsigned(16#2B#, 8);
  gmul3_4(25) <= to_unsigned(16#2E#, 8);
  gmul3_4(26) <= to_unsigned(16#2D#, 8);
  gmul3_4(27) <= to_unsigned(16#24#, 8);
  gmul3_4(28) <= to_unsigned(16#27#, 8);
  gmul3_4(29) <= to_unsigned(16#22#, 8);
  gmul3_4(30) <= to_unsigned(16#21#, 8);
  gmul3_4(31) <= to_unsigned(16#60#, 8);
  gmul3_4(32) <= to_unsigned(16#63#, 8);
  gmul3_4(33) <= to_unsigned(16#66#, 8);
  gmul3_4(34) <= to_unsigned(16#65#, 8);
  gmul3_4(35) <= to_unsigned(16#6C#, 8);
  gmul3_4(36) <= to_unsigned(16#6F#, 8);
  gmul3_4(37) <= to_unsigned(16#6A#, 8);
  gmul3_4(38) <= to_unsigned(16#69#, 8);
  gmul3_4(39) <= to_unsigned(16#78#, 8);
  gmul3_4(40) <= to_unsigned(16#7B#, 8);
  gmul3_4(41) <= to_unsigned(16#7E#, 8);
  gmul3_4(42) <= to_unsigned(16#7D#, 8);
  gmul3_4(43) <= to_unsigned(16#74#, 8);
  gmul3_4(44) <= to_unsigned(16#77#, 8);
  gmul3_4(45) <= to_unsigned(16#72#, 8);
  gmul3_4(46) <= to_unsigned(16#71#, 8);
  gmul3_4(47) <= to_unsigned(16#50#, 8);
  gmul3_4(48) <= to_unsigned(16#53#, 8);
  gmul3_4(49) <= to_unsigned(16#56#, 8);
  gmul3_4(50) <= to_unsigned(16#55#, 8);
  gmul3_4(51) <= to_unsigned(16#5C#, 8);
  gmul3_4(52) <= to_unsigned(16#5F#, 8);
  gmul3_4(53) <= to_unsigned(16#5A#, 8);
  gmul3_4(54) <= to_unsigned(16#59#, 8);
  gmul3_4(55) <= to_unsigned(16#48#, 8);
  gmul3_4(56) <= to_unsigned(16#4B#, 8);
  gmul3_4(57) <= to_unsigned(16#4E#, 8);
  gmul3_4(58) <= to_unsigned(16#4D#, 8);
  gmul3_4(59) <= to_unsigned(16#44#, 8);
  gmul3_4(60) <= to_unsigned(16#47#, 8);
  gmul3_4(61) <= to_unsigned(16#42#, 8);
  gmul3_4(62) <= to_unsigned(16#41#, 8);
  gmul3_4(63) <= to_unsigned(16#C0#, 8);
  gmul3_4(64) <= to_unsigned(16#C3#, 8);
  gmul3_4(65) <= to_unsigned(16#C6#, 8);
  gmul3_4(66) <= to_unsigned(16#C5#, 8);
  gmul3_4(67) <= to_unsigned(16#CC#, 8);
  gmul3_4(68) <= to_unsigned(16#CF#, 8);
  gmul3_4(69) <= to_unsigned(16#CA#, 8);
  gmul3_4(70) <= to_unsigned(16#C9#, 8);
  gmul3_4(71) <= to_unsigned(16#D8#, 8);
  gmul3_4(72) <= to_unsigned(16#DB#, 8);
  gmul3_4(73) <= to_unsigned(16#DE#, 8);
  gmul3_4(74) <= to_unsigned(16#DD#, 8);
  gmul3_4(75) <= to_unsigned(16#D4#, 8);
  gmul3_4(76) <= to_unsigned(16#D7#, 8);
  gmul3_4(77) <= to_unsigned(16#D2#, 8);
  gmul3_4(78) <= to_unsigned(16#D1#, 8);
  gmul3_4(79) <= to_unsigned(16#F0#, 8);
  gmul3_4(80) <= to_unsigned(16#F3#, 8);
  gmul3_4(81) <= to_unsigned(16#F6#, 8);
  gmul3_4(82) <= to_unsigned(16#F5#, 8);
  gmul3_4(83) <= to_unsigned(16#FC#, 8);
  gmul3_4(84) <= to_unsigned(16#FF#, 8);
  gmul3_4(85) <= to_unsigned(16#FA#, 8);
  gmul3_4(86) <= to_unsigned(16#F9#, 8);
  gmul3_4(87) <= to_unsigned(16#E8#, 8);
  gmul3_4(88) <= to_unsigned(16#EB#, 8);
  gmul3_4(89) <= to_unsigned(16#EE#, 8);
  gmul3_4(90) <= to_unsigned(16#ED#, 8);
  gmul3_4(91) <= to_unsigned(16#E4#, 8);
  gmul3_4(92) <= to_unsigned(16#E7#, 8);
  gmul3_4(93) <= to_unsigned(16#E2#, 8);
  gmul3_4(94) <= to_unsigned(16#E1#, 8);
  gmul3_4(95) <= to_unsigned(16#A0#, 8);
  gmul3_4(96) <= to_unsigned(16#A3#, 8);
  gmul3_4(97) <= to_unsigned(16#A6#, 8);
  gmul3_4(98) <= to_unsigned(16#A5#, 8);
  gmul3_4(99) <= to_unsigned(16#AC#, 8);
  gmul3_4(100) <= to_unsigned(16#AF#, 8);
  gmul3_4(101) <= to_unsigned(16#AA#, 8);
  gmul3_4(102) <= to_unsigned(16#A9#, 8);
  gmul3_4(103) <= to_unsigned(16#B8#, 8);
  gmul3_4(104) <= to_unsigned(16#BB#, 8);
  gmul3_4(105) <= to_unsigned(16#BE#, 8);
  gmul3_4(106) <= to_unsigned(16#BD#, 8);
  gmul3_4(107) <= to_unsigned(16#B4#, 8);
  gmul3_4(108) <= to_unsigned(16#B7#, 8);
  gmul3_4(109) <= to_unsigned(16#B2#, 8);
  gmul3_4(110) <= to_unsigned(16#B1#, 8);
  gmul3_4(111) <= to_unsigned(16#90#, 8);
  gmul3_4(112) <= to_unsigned(16#93#, 8);
  gmul3_4(113) <= to_unsigned(16#96#, 8);
  gmul3_4(114) <= to_unsigned(16#95#, 8);
  gmul3_4(115) <= to_unsigned(16#9C#, 8);
  gmul3_4(116) <= to_unsigned(16#9F#, 8);
  gmul3_4(117) <= to_unsigned(16#9A#, 8);
  gmul3_4(118) <= to_unsigned(16#99#, 8);
  gmul3_4(119) <= to_unsigned(16#88#, 8);
  gmul3_4(120) <= to_unsigned(16#8B#, 8);
  gmul3_4(121) <= to_unsigned(16#8E#, 8);
  gmul3_4(122) <= to_unsigned(16#8D#, 8);
  gmul3_4(123) <= to_unsigned(16#84#, 8);
  gmul3_4(124) <= to_unsigned(16#87#, 8);
  gmul3_4(125) <= to_unsigned(16#82#, 8);
  gmul3_4(126) <= to_unsigned(16#81#, 8);
  gmul3_4(127) <= to_unsigned(16#9B#, 8);
  gmul3_4(128) <= to_unsigned(16#98#, 8);
  gmul3_4(129) <= to_unsigned(16#9D#, 8);
  gmul3_4(130) <= to_unsigned(16#9E#, 8);
  gmul3_4(131) <= to_unsigned(16#97#, 8);
  gmul3_4(132) <= to_unsigned(16#94#, 8);
  gmul3_4(133) <= to_unsigned(16#91#, 8);
  gmul3_4(134) <= to_unsigned(16#92#, 8);
  gmul3_4(135) <= to_unsigned(16#83#, 8);
  gmul3_4(136) <= to_unsigned(16#80#, 8);
  gmul3_4(137) <= to_unsigned(16#85#, 8);
  gmul3_4(138) <= to_unsigned(16#86#, 8);
  gmul3_4(139) <= to_unsigned(16#8F#, 8);
  gmul3_4(140) <= to_unsigned(16#8C#, 8);
  gmul3_4(141) <= to_unsigned(16#89#, 8);
  gmul3_4(142) <= to_unsigned(16#8A#, 8);
  gmul3_4(143) <= to_unsigned(16#AB#, 8);
  gmul3_4(144) <= to_unsigned(16#A8#, 8);
  gmul3_4(145) <= to_unsigned(16#AD#, 8);
  gmul3_4(146) <= to_unsigned(16#AE#, 8);
  gmul3_4(147) <= to_unsigned(16#A7#, 8);
  gmul3_4(148) <= to_unsigned(16#A4#, 8);
  gmul3_4(149) <= to_unsigned(16#A1#, 8);
  gmul3_4(150) <= to_unsigned(16#A2#, 8);
  gmul3_4(151) <= to_unsigned(16#B3#, 8);
  gmul3_4(152) <= to_unsigned(16#B0#, 8);
  gmul3_4(153) <= to_unsigned(16#B5#, 8);
  gmul3_4(154) <= to_unsigned(16#B6#, 8);
  gmul3_4(155) <= to_unsigned(16#BF#, 8);
  gmul3_4(156) <= to_unsigned(16#BC#, 8);
  gmul3_4(157) <= to_unsigned(16#B9#, 8);
  gmul3_4(158) <= to_unsigned(16#BA#, 8);
  gmul3_4(159) <= to_unsigned(16#FB#, 8);
  gmul3_4(160) <= to_unsigned(16#F8#, 8);
  gmul3_4(161) <= to_unsigned(16#FD#, 8);
  gmul3_4(162) <= to_unsigned(16#FE#, 8);
  gmul3_4(163) <= to_unsigned(16#F7#, 8);
  gmul3_4(164) <= to_unsigned(16#F4#, 8);
  gmul3_4(165) <= to_unsigned(16#F1#, 8);
  gmul3_4(166) <= to_unsigned(16#F2#, 8);
  gmul3_4(167) <= to_unsigned(16#E3#, 8);
  gmul3_4(168) <= to_unsigned(16#E0#, 8);
  gmul3_4(169) <= to_unsigned(16#E5#, 8);
  gmul3_4(170) <= to_unsigned(16#E6#, 8);
  gmul3_4(171) <= to_unsigned(16#EF#, 8);
  gmul3_4(172) <= to_unsigned(16#EC#, 8);
  gmul3_4(173) <= to_unsigned(16#E9#, 8);
  gmul3_4(174) <= to_unsigned(16#EA#, 8);
  gmul3_4(175) <= to_unsigned(16#CB#, 8);
  gmul3_4(176) <= to_unsigned(16#C8#, 8);
  gmul3_4(177) <= to_unsigned(16#CD#, 8);
  gmul3_4(178) <= to_unsigned(16#CE#, 8);
  gmul3_4(179) <= to_unsigned(16#C7#, 8);
  gmul3_4(180) <= to_unsigned(16#C4#, 8);
  gmul3_4(181) <= to_unsigned(16#C1#, 8);
  gmul3_4(182) <= to_unsigned(16#C2#, 8);
  gmul3_4(183) <= to_unsigned(16#D3#, 8);
  gmul3_4(184) <= to_unsigned(16#D0#, 8);
  gmul3_4(185) <= to_unsigned(16#D5#, 8);
  gmul3_4(186) <= to_unsigned(16#D6#, 8);
  gmul3_4(187) <= to_unsigned(16#DF#, 8);
  gmul3_4(188) <= to_unsigned(16#DC#, 8);
  gmul3_4(189) <= to_unsigned(16#D9#, 8);
  gmul3_4(190) <= to_unsigned(16#DA#, 8);
  gmul3_4(191) <= to_unsigned(16#5B#, 8);
  gmul3_4(192) <= to_unsigned(16#58#, 8);
  gmul3_4(193) <= to_unsigned(16#5D#, 8);
  gmul3_4(194) <= to_unsigned(16#5E#, 8);
  gmul3_4(195) <= to_unsigned(16#57#, 8);
  gmul3_4(196) <= to_unsigned(16#54#, 8);
  gmul3_4(197) <= to_unsigned(16#51#, 8);
  gmul3_4(198) <= to_unsigned(16#52#, 8);
  gmul3_4(199) <= to_unsigned(16#43#, 8);
  gmul3_4(200) <= to_unsigned(16#40#, 8);
  gmul3_4(201) <= to_unsigned(16#45#, 8);
  gmul3_4(202) <= to_unsigned(16#46#, 8);
  gmul3_4(203) <= to_unsigned(16#4F#, 8);
  gmul3_4(204) <= to_unsigned(16#4C#, 8);
  gmul3_4(205) <= to_unsigned(16#49#, 8);
  gmul3_4(206) <= to_unsigned(16#4A#, 8);
  gmul3_4(207) <= to_unsigned(16#6B#, 8);
  gmul3_4(208) <= to_unsigned(16#68#, 8);
  gmul3_4(209) <= to_unsigned(16#6D#, 8);
  gmul3_4(210) <= to_unsigned(16#6E#, 8);
  gmul3_4(211) <= to_unsigned(16#67#, 8);
  gmul3_4(212) <= to_unsigned(16#64#, 8);
  gmul3_4(213) <= to_unsigned(16#61#, 8);
  gmul3_4(214) <= to_unsigned(16#62#, 8);
  gmul3_4(215) <= to_unsigned(16#73#, 8);
  gmul3_4(216) <= to_unsigned(16#70#, 8);
  gmul3_4(217) <= to_unsigned(16#75#, 8);
  gmul3_4(218) <= to_unsigned(16#76#, 8);
  gmul3_4(219) <= to_unsigned(16#7F#, 8);
  gmul3_4(220) <= to_unsigned(16#7C#, 8);
  gmul3_4(221) <= to_unsigned(16#79#, 8);
  gmul3_4(222) <= to_unsigned(16#7A#, 8);
  gmul3_4(223) <= to_unsigned(16#3B#, 8);
  gmul3_4(224) <= to_unsigned(16#38#, 8);
  gmul3_4(225) <= to_unsigned(16#3D#, 8);
  gmul3_4(226) <= to_unsigned(16#3E#, 8);
  gmul3_4(227) <= to_unsigned(16#37#, 8);
  gmul3_4(228) <= to_unsigned(16#34#, 8);
  gmul3_4(229) <= to_unsigned(16#31#, 8);
  gmul3_4(230) <= to_unsigned(16#32#, 8);
  gmul3_4(231) <= to_unsigned(16#23#, 8);
  gmul3_4(232) <= to_unsigned(16#20#, 8);
  gmul3_4(233) <= to_unsigned(16#25#, 8);
  gmul3_4(234) <= to_unsigned(16#26#, 8);
  gmul3_4(235) <= to_unsigned(16#2F#, 8);
  gmul3_4(236) <= to_unsigned(16#2C#, 8);
  gmul3_4(237) <= to_unsigned(16#29#, 8);
  gmul3_4(238) <= to_unsigned(16#2A#, 8);
  gmul3_4(239) <= to_unsigned(16#0B#, 8);
  gmul3_4(240) <= to_unsigned(16#08#, 8);
  gmul3_4(241) <= to_unsigned(16#0D#, 8);
  gmul3_4(242) <= to_unsigned(16#0E#, 8);
  gmul3_4(243) <= to_unsigned(16#07#, 8);
  gmul3_4(244) <= to_unsigned(16#04#, 8);
  gmul3_4(245) <= to_unsigned(16#01#, 8);
  gmul3_4(246) <= to_unsigned(16#02#, 8);
  gmul3_4(247) <= to_unsigned(16#13#, 8);
  gmul3_4(248) <= to_unsigned(16#10#, 8);
  gmul3_4(249) <= to_unsigned(16#15#, 8);
  gmul3_4(250) <= to_unsigned(16#16#, 8);
  gmul3_4(251) <= to_unsigned(16#1F#, 8);
  gmul3_4(252) <= to_unsigned(16#1C#, 8);
  gmul3_4(253) <= to_unsigned(16#19#, 8);
  gmul3_4(254) <= to_unsigned(16#1A#, 8);
  gmul3_4(255) <= to_unsigned(16#1A#, 8);

  gmul2_5(0) <= to_unsigned(16#02#, 8);
  gmul2_5(1) <= to_unsigned(16#04#, 8);
  gmul2_5(2) <= to_unsigned(16#06#, 8);
  gmul2_5(3) <= to_unsigned(16#08#, 8);
  gmul2_5(4) <= to_unsigned(16#0A#, 8);
  gmul2_5(5) <= to_unsigned(16#0C#, 8);
  gmul2_5(6) <= to_unsigned(16#0E#, 8);
  gmul2_5(7) <= to_unsigned(16#10#, 8);
  gmul2_5(8) <= to_unsigned(16#12#, 8);
  gmul2_5(9) <= to_unsigned(16#14#, 8);
  gmul2_5(10) <= to_unsigned(16#16#, 8);
  gmul2_5(11) <= to_unsigned(16#18#, 8);
  gmul2_5(12) <= to_unsigned(16#1A#, 8);
  gmul2_5(13) <= to_unsigned(16#1C#, 8);
  gmul2_5(14) <= to_unsigned(16#1E#, 8);
  gmul2_5(15) <= to_unsigned(16#20#, 8);
  gmul2_5(16) <= to_unsigned(16#22#, 8);
  gmul2_5(17) <= to_unsigned(16#24#, 8);
  gmul2_5(18) <= to_unsigned(16#26#, 8);
  gmul2_5(19) <= to_unsigned(16#28#, 8);
  gmul2_5(20) <= to_unsigned(16#2A#, 8);
  gmul2_5(21) <= to_unsigned(16#2C#, 8);
  gmul2_5(22) <= to_unsigned(16#2E#, 8);
  gmul2_5(23) <= to_unsigned(16#30#, 8);
  gmul2_5(24) <= to_unsigned(16#32#, 8);
  gmul2_5(25) <= to_unsigned(16#34#, 8);
  gmul2_5(26) <= to_unsigned(16#36#, 8);
  gmul2_5(27) <= to_unsigned(16#38#, 8);
  gmul2_5(28) <= to_unsigned(16#3A#, 8);
  gmul2_5(29) <= to_unsigned(16#3C#, 8);
  gmul2_5(30) <= to_unsigned(16#3E#, 8);
  gmul2_5(31) <= to_unsigned(16#40#, 8);
  gmul2_5(32) <= to_unsigned(16#42#, 8);
  gmul2_5(33) <= to_unsigned(16#44#, 8);
  gmul2_5(34) <= to_unsigned(16#46#, 8);
  gmul2_5(35) <= to_unsigned(16#48#, 8);
  gmul2_5(36) <= to_unsigned(16#4A#, 8);
  gmul2_5(37) <= to_unsigned(16#4C#, 8);
  gmul2_5(38) <= to_unsigned(16#4E#, 8);
  gmul2_5(39) <= to_unsigned(16#50#, 8);
  gmul2_5(40) <= to_unsigned(16#52#, 8);
  gmul2_5(41) <= to_unsigned(16#54#, 8);
  gmul2_5(42) <= to_unsigned(16#56#, 8);
  gmul2_5(43) <= to_unsigned(16#58#, 8);
  gmul2_5(44) <= to_unsigned(16#5A#, 8);
  gmul2_5(45) <= to_unsigned(16#5C#, 8);
  gmul2_5(46) <= to_unsigned(16#5E#, 8);
  gmul2_5(47) <= to_unsigned(16#60#, 8);
  gmul2_5(48) <= to_unsigned(16#62#, 8);
  gmul2_5(49) <= to_unsigned(16#64#, 8);
  gmul2_5(50) <= to_unsigned(16#66#, 8);
  gmul2_5(51) <= to_unsigned(16#68#, 8);
  gmul2_5(52) <= to_unsigned(16#6A#, 8);
  gmul2_5(53) <= to_unsigned(16#6C#, 8);
  gmul2_5(54) <= to_unsigned(16#6E#, 8);
  gmul2_5(55) <= to_unsigned(16#70#, 8);
  gmul2_5(56) <= to_unsigned(16#72#, 8);
  gmul2_5(57) <= to_unsigned(16#74#, 8);
  gmul2_5(58) <= to_unsigned(16#76#, 8);
  gmul2_5(59) <= to_unsigned(16#78#, 8);
  gmul2_5(60) <= to_unsigned(16#7A#, 8);
  gmul2_5(61) <= to_unsigned(16#7C#, 8);
  gmul2_5(62) <= to_unsigned(16#7E#, 8);
  gmul2_5(63) <= to_unsigned(16#80#, 8);
  gmul2_5(64) <= to_unsigned(16#82#, 8);
  gmul2_5(65) <= to_unsigned(16#84#, 8);
  gmul2_5(66) <= to_unsigned(16#86#, 8);
  gmul2_5(67) <= to_unsigned(16#88#, 8);
  gmul2_5(68) <= to_unsigned(16#8A#, 8);
  gmul2_5(69) <= to_unsigned(16#8C#, 8);
  gmul2_5(70) <= to_unsigned(16#8E#, 8);
  gmul2_5(71) <= to_unsigned(16#90#, 8);
  gmul2_5(72) <= to_unsigned(16#92#, 8);
  gmul2_5(73) <= to_unsigned(16#94#, 8);
  gmul2_5(74) <= to_unsigned(16#96#, 8);
  gmul2_5(75) <= to_unsigned(16#98#, 8);
  gmul2_5(76) <= to_unsigned(16#9A#, 8);
  gmul2_5(77) <= to_unsigned(16#9C#, 8);
  gmul2_5(78) <= to_unsigned(16#9E#, 8);
  gmul2_5(79) <= to_unsigned(16#A0#, 8);
  gmul2_5(80) <= to_unsigned(16#A2#, 8);
  gmul2_5(81) <= to_unsigned(16#A4#, 8);
  gmul2_5(82) <= to_unsigned(16#A6#, 8);
  gmul2_5(83) <= to_unsigned(16#A8#, 8);
  gmul2_5(84) <= to_unsigned(16#AA#, 8);
  gmul2_5(85) <= to_unsigned(16#AC#, 8);
  gmul2_5(86) <= to_unsigned(16#AE#, 8);
  gmul2_5(87) <= to_unsigned(16#B0#, 8);
  gmul2_5(88) <= to_unsigned(16#B2#, 8);
  gmul2_5(89) <= to_unsigned(16#B4#, 8);
  gmul2_5(90) <= to_unsigned(16#B6#, 8);
  gmul2_5(91) <= to_unsigned(16#B8#, 8);
  gmul2_5(92) <= to_unsigned(16#BA#, 8);
  gmul2_5(93) <= to_unsigned(16#BC#, 8);
  gmul2_5(94) <= to_unsigned(16#BE#, 8);
  gmul2_5(95) <= to_unsigned(16#C0#, 8);
  gmul2_5(96) <= to_unsigned(16#C2#, 8);
  gmul2_5(97) <= to_unsigned(16#C4#, 8);
  gmul2_5(98) <= to_unsigned(16#C6#, 8);
  gmul2_5(99) <= to_unsigned(16#C8#, 8);
  gmul2_5(100) <= to_unsigned(16#CA#, 8);
  gmul2_5(101) <= to_unsigned(16#CC#, 8);
  gmul2_5(102) <= to_unsigned(16#CE#, 8);
  gmul2_5(103) <= to_unsigned(16#D0#, 8);
  gmul2_5(104) <= to_unsigned(16#D2#, 8);
  gmul2_5(105) <= to_unsigned(16#D4#, 8);
  gmul2_5(106) <= to_unsigned(16#D6#, 8);
  gmul2_5(107) <= to_unsigned(16#D8#, 8);
  gmul2_5(108) <= to_unsigned(16#DA#, 8);
  gmul2_5(109) <= to_unsigned(16#DC#, 8);
  gmul2_5(110) <= to_unsigned(16#DE#, 8);
  gmul2_5(111) <= to_unsigned(16#E0#, 8);
  gmul2_5(112) <= to_unsigned(16#E2#, 8);
  gmul2_5(113) <= to_unsigned(16#E4#, 8);
  gmul2_5(114) <= to_unsigned(16#E6#, 8);
  gmul2_5(115) <= to_unsigned(16#E8#, 8);
  gmul2_5(116) <= to_unsigned(16#EA#, 8);
  gmul2_5(117) <= to_unsigned(16#EC#, 8);
  gmul2_5(118) <= to_unsigned(16#EE#, 8);
  gmul2_5(119) <= to_unsigned(16#F0#, 8);
  gmul2_5(120) <= to_unsigned(16#F2#, 8);
  gmul2_5(121) <= to_unsigned(16#F4#, 8);
  gmul2_5(122) <= to_unsigned(16#F6#, 8);
  gmul2_5(123) <= to_unsigned(16#F8#, 8);
  gmul2_5(124) <= to_unsigned(16#FA#, 8);
  gmul2_5(125) <= to_unsigned(16#FC#, 8);
  gmul2_5(126) <= to_unsigned(16#FE#, 8);
  gmul2_5(127) <= to_unsigned(16#1B#, 8);
  gmul2_5(128) <= to_unsigned(16#19#, 8);
  gmul2_5(129) <= to_unsigned(16#1F#, 8);
  gmul2_5(130) <= to_unsigned(16#1D#, 8);
  gmul2_5(131) <= to_unsigned(16#13#, 8);
  gmul2_5(132) <= to_unsigned(16#11#, 8);
  gmul2_5(133) <= to_unsigned(16#17#, 8);
  gmul2_5(134) <= to_unsigned(16#15#, 8);
  gmul2_5(135) <= to_unsigned(16#0B#, 8);
  gmul2_5(136) <= to_unsigned(16#09#, 8);
  gmul2_5(137) <= to_unsigned(16#0F#, 8);
  gmul2_5(138) <= to_unsigned(16#0D#, 8);
  gmul2_5(139) <= to_unsigned(16#03#, 8);
  gmul2_5(140) <= to_unsigned(16#01#, 8);
  gmul2_5(141) <= to_unsigned(16#07#, 8);
  gmul2_5(142) <= to_unsigned(16#05#, 8);
  gmul2_5(143) <= to_unsigned(16#3B#, 8);
  gmul2_5(144) <= to_unsigned(16#39#, 8);
  gmul2_5(145) <= to_unsigned(16#3F#, 8);
  gmul2_5(146) <= to_unsigned(16#3D#, 8);
  gmul2_5(147) <= to_unsigned(16#33#, 8);
  gmul2_5(148) <= to_unsigned(16#31#, 8);
  gmul2_5(149) <= to_unsigned(16#37#, 8);
  gmul2_5(150) <= to_unsigned(16#35#, 8);
  gmul2_5(151) <= to_unsigned(16#2B#, 8);
  gmul2_5(152) <= to_unsigned(16#29#, 8);
  gmul2_5(153) <= to_unsigned(16#2F#, 8);
  gmul2_5(154) <= to_unsigned(16#2D#, 8);
  gmul2_5(155) <= to_unsigned(16#23#, 8);
  gmul2_5(156) <= to_unsigned(16#21#, 8);
  gmul2_5(157) <= to_unsigned(16#27#, 8);
  gmul2_5(158) <= to_unsigned(16#25#, 8);
  gmul2_5(159) <= to_unsigned(16#5B#, 8);
  gmul2_5(160) <= to_unsigned(16#59#, 8);
  gmul2_5(161) <= to_unsigned(16#5F#, 8);
  gmul2_5(162) <= to_unsigned(16#5D#, 8);
  gmul2_5(163) <= to_unsigned(16#53#, 8);
  gmul2_5(164) <= to_unsigned(16#51#, 8);
  gmul2_5(165) <= to_unsigned(16#57#, 8);
  gmul2_5(166) <= to_unsigned(16#55#, 8);
  gmul2_5(167) <= to_unsigned(16#4B#, 8);
  gmul2_5(168) <= to_unsigned(16#49#, 8);
  gmul2_5(169) <= to_unsigned(16#4F#, 8);
  gmul2_5(170) <= to_unsigned(16#4D#, 8);
  gmul2_5(171) <= to_unsigned(16#43#, 8);
  gmul2_5(172) <= to_unsigned(16#41#, 8);
  gmul2_5(173) <= to_unsigned(16#47#, 8);
  gmul2_5(174) <= to_unsigned(16#45#, 8);
  gmul2_5(175) <= to_unsigned(16#7B#, 8);
  gmul2_5(176) <= to_unsigned(16#79#, 8);
  gmul2_5(177) <= to_unsigned(16#7F#, 8);
  gmul2_5(178) <= to_unsigned(16#7D#, 8);
  gmul2_5(179) <= to_unsigned(16#73#, 8);
  gmul2_5(180) <= to_unsigned(16#71#, 8);
  gmul2_5(181) <= to_unsigned(16#77#, 8);
  gmul2_5(182) <= to_unsigned(16#75#, 8);
  gmul2_5(183) <= to_unsigned(16#6B#, 8);
  gmul2_5(184) <= to_unsigned(16#69#, 8);
  gmul2_5(185) <= to_unsigned(16#6F#, 8);
  gmul2_5(186) <= to_unsigned(16#6D#, 8);
  gmul2_5(187) <= to_unsigned(16#63#, 8);
  gmul2_5(188) <= to_unsigned(16#61#, 8);
  gmul2_5(189) <= to_unsigned(16#67#, 8);
  gmul2_5(190) <= to_unsigned(16#65#, 8);
  gmul2_5(191) <= to_unsigned(16#9B#, 8);
  gmul2_5(192) <= to_unsigned(16#99#, 8);
  gmul2_5(193) <= to_unsigned(16#9F#, 8);
  gmul2_5(194) <= to_unsigned(16#9D#, 8);
  gmul2_5(195) <= to_unsigned(16#93#, 8);
  gmul2_5(196) <= to_unsigned(16#91#, 8);
  gmul2_5(197) <= to_unsigned(16#97#, 8);
  gmul2_5(198) <= to_unsigned(16#95#, 8);
  gmul2_5(199) <= to_unsigned(16#8B#, 8);
  gmul2_5(200) <= to_unsigned(16#89#, 8);
  gmul2_5(201) <= to_unsigned(16#8F#, 8);
  gmul2_5(202) <= to_unsigned(16#8D#, 8);
  gmul2_5(203) <= to_unsigned(16#83#, 8);
  gmul2_5(204) <= to_unsigned(16#81#, 8);
  gmul2_5(205) <= to_unsigned(16#87#, 8);
  gmul2_5(206) <= to_unsigned(16#85#, 8);
  gmul2_5(207) <= to_unsigned(16#BB#, 8);
  gmul2_5(208) <= to_unsigned(16#B9#, 8);
  gmul2_5(209) <= to_unsigned(16#BF#, 8);
  gmul2_5(210) <= to_unsigned(16#BD#, 8);
  gmul2_5(211) <= to_unsigned(16#B3#, 8);
  gmul2_5(212) <= to_unsigned(16#B1#, 8);
  gmul2_5(213) <= to_unsigned(16#B7#, 8);
  gmul2_5(214) <= to_unsigned(16#B5#, 8);
  gmul2_5(215) <= to_unsigned(16#AB#, 8);
  gmul2_5(216) <= to_unsigned(16#A9#, 8);
  gmul2_5(217) <= to_unsigned(16#AF#, 8);
  gmul2_5(218) <= to_unsigned(16#AD#, 8);
  gmul2_5(219) <= to_unsigned(16#A3#, 8);
  gmul2_5(220) <= to_unsigned(16#A1#, 8);
  gmul2_5(221) <= to_unsigned(16#A7#, 8);
  gmul2_5(222) <= to_unsigned(16#A5#, 8);
  gmul2_5(223) <= to_unsigned(16#DB#, 8);
  gmul2_5(224) <= to_unsigned(16#D9#, 8);
  gmul2_5(225) <= to_unsigned(16#DF#, 8);
  gmul2_5(226) <= to_unsigned(16#DD#, 8);
  gmul2_5(227) <= to_unsigned(16#D3#, 8);
  gmul2_5(228) <= to_unsigned(16#D1#, 8);
  gmul2_5(229) <= to_unsigned(16#D7#, 8);
  gmul2_5(230) <= to_unsigned(16#D5#, 8);
  gmul2_5(231) <= to_unsigned(16#CB#, 8);
  gmul2_5(232) <= to_unsigned(16#C9#, 8);
  gmul2_5(233) <= to_unsigned(16#CF#, 8);
  gmul2_5(234) <= to_unsigned(16#CD#, 8);
  gmul2_5(235) <= to_unsigned(16#C3#, 8);
  gmul2_5(236) <= to_unsigned(16#C1#, 8);
  gmul2_5(237) <= to_unsigned(16#C7#, 8);
  gmul2_5(238) <= to_unsigned(16#C5#, 8);
  gmul2_5(239) <= to_unsigned(16#FB#, 8);
  gmul2_5(240) <= to_unsigned(16#F9#, 8);
  gmul2_5(241) <= to_unsigned(16#FF#, 8);
  gmul2_5(242) <= to_unsigned(16#FD#, 8);
  gmul2_5(243) <= to_unsigned(16#F3#, 8);
  gmul2_5(244) <= to_unsigned(16#F1#, 8);
  gmul2_5(245) <= to_unsigned(16#F7#, 8);
  gmul2_5(246) <= to_unsigned(16#F5#, 8);
  gmul2_5(247) <= to_unsigned(16#EB#, 8);
  gmul2_5(248) <= to_unsigned(16#E9#, 8);
  gmul2_5(249) <= to_unsigned(16#EF#, 8);
  gmul2_5(250) <= to_unsigned(16#ED#, 8);
  gmul2_5(251) <= to_unsigned(16#E3#, 8);
  gmul2_5(252) <= to_unsigned(16#E1#, 8);
  gmul2_5(253) <= to_unsigned(16#E7#, 8);
  gmul2_5(254) <= to_unsigned(16#E5#, 8);
  gmul2_5(255) <= to_unsigned(16#E5#, 8);

  gmul3_5(0) <= to_unsigned(16#03#, 8);
  gmul3_5(1) <= to_unsigned(16#06#, 8);
  gmul3_5(2) <= to_unsigned(16#05#, 8);
  gmul3_5(3) <= to_unsigned(16#0C#, 8);
  gmul3_5(4) <= to_unsigned(16#0F#, 8);
  gmul3_5(5) <= to_unsigned(16#0A#, 8);
  gmul3_5(6) <= to_unsigned(16#09#, 8);
  gmul3_5(7) <= to_unsigned(16#18#, 8);
  gmul3_5(8) <= to_unsigned(16#1B#, 8);
  gmul3_5(9) <= to_unsigned(16#1E#, 8);
  gmul3_5(10) <= to_unsigned(16#1D#, 8);
  gmul3_5(11) <= to_unsigned(16#14#, 8);
  gmul3_5(12) <= to_unsigned(16#17#, 8);
  gmul3_5(13) <= to_unsigned(16#12#, 8);
  gmul3_5(14) <= to_unsigned(16#11#, 8);
  gmul3_5(15) <= to_unsigned(16#30#, 8);
  gmul3_5(16) <= to_unsigned(16#33#, 8);
  gmul3_5(17) <= to_unsigned(16#36#, 8);
  gmul3_5(18) <= to_unsigned(16#35#, 8);
  gmul3_5(19) <= to_unsigned(16#3C#, 8);
  gmul3_5(20) <= to_unsigned(16#3F#, 8);
  gmul3_5(21) <= to_unsigned(16#3A#, 8);
  gmul3_5(22) <= to_unsigned(16#39#, 8);
  gmul3_5(23) <= to_unsigned(16#28#, 8);
  gmul3_5(24) <= to_unsigned(16#2B#, 8);
  gmul3_5(25) <= to_unsigned(16#2E#, 8);
  gmul3_5(26) <= to_unsigned(16#2D#, 8);
  gmul3_5(27) <= to_unsigned(16#24#, 8);
  gmul3_5(28) <= to_unsigned(16#27#, 8);
  gmul3_5(29) <= to_unsigned(16#22#, 8);
  gmul3_5(30) <= to_unsigned(16#21#, 8);
  gmul3_5(31) <= to_unsigned(16#60#, 8);
  gmul3_5(32) <= to_unsigned(16#63#, 8);
  gmul3_5(33) <= to_unsigned(16#66#, 8);
  gmul3_5(34) <= to_unsigned(16#65#, 8);
  gmul3_5(35) <= to_unsigned(16#6C#, 8);
  gmul3_5(36) <= to_unsigned(16#6F#, 8);
  gmul3_5(37) <= to_unsigned(16#6A#, 8);
  gmul3_5(38) <= to_unsigned(16#69#, 8);
  gmul3_5(39) <= to_unsigned(16#78#, 8);
  gmul3_5(40) <= to_unsigned(16#7B#, 8);
  gmul3_5(41) <= to_unsigned(16#7E#, 8);
  gmul3_5(42) <= to_unsigned(16#7D#, 8);
  gmul3_5(43) <= to_unsigned(16#74#, 8);
  gmul3_5(44) <= to_unsigned(16#77#, 8);
  gmul3_5(45) <= to_unsigned(16#72#, 8);
  gmul3_5(46) <= to_unsigned(16#71#, 8);
  gmul3_5(47) <= to_unsigned(16#50#, 8);
  gmul3_5(48) <= to_unsigned(16#53#, 8);
  gmul3_5(49) <= to_unsigned(16#56#, 8);
  gmul3_5(50) <= to_unsigned(16#55#, 8);
  gmul3_5(51) <= to_unsigned(16#5C#, 8);
  gmul3_5(52) <= to_unsigned(16#5F#, 8);
  gmul3_5(53) <= to_unsigned(16#5A#, 8);
  gmul3_5(54) <= to_unsigned(16#59#, 8);
  gmul3_5(55) <= to_unsigned(16#48#, 8);
  gmul3_5(56) <= to_unsigned(16#4B#, 8);
  gmul3_5(57) <= to_unsigned(16#4E#, 8);
  gmul3_5(58) <= to_unsigned(16#4D#, 8);
  gmul3_5(59) <= to_unsigned(16#44#, 8);
  gmul3_5(60) <= to_unsigned(16#47#, 8);
  gmul3_5(61) <= to_unsigned(16#42#, 8);
  gmul3_5(62) <= to_unsigned(16#41#, 8);
  gmul3_5(63) <= to_unsigned(16#C0#, 8);
  gmul3_5(64) <= to_unsigned(16#C3#, 8);
  gmul3_5(65) <= to_unsigned(16#C6#, 8);
  gmul3_5(66) <= to_unsigned(16#C5#, 8);
  gmul3_5(67) <= to_unsigned(16#CC#, 8);
  gmul3_5(68) <= to_unsigned(16#CF#, 8);
  gmul3_5(69) <= to_unsigned(16#CA#, 8);
  gmul3_5(70) <= to_unsigned(16#C9#, 8);
  gmul3_5(71) <= to_unsigned(16#D8#, 8);
  gmul3_5(72) <= to_unsigned(16#DB#, 8);
  gmul3_5(73) <= to_unsigned(16#DE#, 8);
  gmul3_5(74) <= to_unsigned(16#DD#, 8);
  gmul3_5(75) <= to_unsigned(16#D4#, 8);
  gmul3_5(76) <= to_unsigned(16#D7#, 8);
  gmul3_5(77) <= to_unsigned(16#D2#, 8);
  gmul3_5(78) <= to_unsigned(16#D1#, 8);
  gmul3_5(79) <= to_unsigned(16#F0#, 8);
  gmul3_5(80) <= to_unsigned(16#F3#, 8);
  gmul3_5(81) <= to_unsigned(16#F6#, 8);
  gmul3_5(82) <= to_unsigned(16#F5#, 8);
  gmul3_5(83) <= to_unsigned(16#FC#, 8);
  gmul3_5(84) <= to_unsigned(16#FF#, 8);
  gmul3_5(85) <= to_unsigned(16#FA#, 8);
  gmul3_5(86) <= to_unsigned(16#F9#, 8);
  gmul3_5(87) <= to_unsigned(16#E8#, 8);
  gmul3_5(88) <= to_unsigned(16#EB#, 8);
  gmul3_5(89) <= to_unsigned(16#EE#, 8);
  gmul3_5(90) <= to_unsigned(16#ED#, 8);
  gmul3_5(91) <= to_unsigned(16#E4#, 8);
  gmul3_5(92) <= to_unsigned(16#E7#, 8);
  gmul3_5(93) <= to_unsigned(16#E2#, 8);
  gmul3_5(94) <= to_unsigned(16#E1#, 8);
  gmul3_5(95) <= to_unsigned(16#A0#, 8);
  gmul3_5(96) <= to_unsigned(16#A3#, 8);
  gmul3_5(97) <= to_unsigned(16#A6#, 8);
  gmul3_5(98) <= to_unsigned(16#A5#, 8);
  gmul3_5(99) <= to_unsigned(16#AC#, 8);
  gmul3_5(100) <= to_unsigned(16#AF#, 8);
  gmul3_5(101) <= to_unsigned(16#AA#, 8);
  gmul3_5(102) <= to_unsigned(16#A9#, 8);
  gmul3_5(103) <= to_unsigned(16#B8#, 8);
  gmul3_5(104) <= to_unsigned(16#BB#, 8);
  gmul3_5(105) <= to_unsigned(16#BE#, 8);
  gmul3_5(106) <= to_unsigned(16#BD#, 8);
  gmul3_5(107) <= to_unsigned(16#B4#, 8);
  gmul3_5(108) <= to_unsigned(16#B7#, 8);
  gmul3_5(109) <= to_unsigned(16#B2#, 8);
  gmul3_5(110) <= to_unsigned(16#B1#, 8);
  gmul3_5(111) <= to_unsigned(16#90#, 8);
  gmul3_5(112) <= to_unsigned(16#93#, 8);
  gmul3_5(113) <= to_unsigned(16#96#, 8);
  gmul3_5(114) <= to_unsigned(16#95#, 8);
  gmul3_5(115) <= to_unsigned(16#9C#, 8);
  gmul3_5(116) <= to_unsigned(16#9F#, 8);
  gmul3_5(117) <= to_unsigned(16#9A#, 8);
  gmul3_5(118) <= to_unsigned(16#99#, 8);
  gmul3_5(119) <= to_unsigned(16#88#, 8);
  gmul3_5(120) <= to_unsigned(16#8B#, 8);
  gmul3_5(121) <= to_unsigned(16#8E#, 8);
  gmul3_5(122) <= to_unsigned(16#8D#, 8);
  gmul3_5(123) <= to_unsigned(16#84#, 8);
  gmul3_5(124) <= to_unsigned(16#87#, 8);
  gmul3_5(125) <= to_unsigned(16#82#, 8);
  gmul3_5(126) <= to_unsigned(16#81#, 8);
  gmul3_5(127) <= to_unsigned(16#9B#, 8);
  gmul3_5(128) <= to_unsigned(16#98#, 8);
  gmul3_5(129) <= to_unsigned(16#9D#, 8);
  gmul3_5(130) <= to_unsigned(16#9E#, 8);
  gmul3_5(131) <= to_unsigned(16#97#, 8);
  gmul3_5(132) <= to_unsigned(16#94#, 8);
  gmul3_5(133) <= to_unsigned(16#91#, 8);
  gmul3_5(134) <= to_unsigned(16#92#, 8);
  gmul3_5(135) <= to_unsigned(16#83#, 8);
  gmul3_5(136) <= to_unsigned(16#80#, 8);
  gmul3_5(137) <= to_unsigned(16#85#, 8);
  gmul3_5(138) <= to_unsigned(16#86#, 8);
  gmul3_5(139) <= to_unsigned(16#8F#, 8);
  gmul3_5(140) <= to_unsigned(16#8C#, 8);
  gmul3_5(141) <= to_unsigned(16#89#, 8);
  gmul3_5(142) <= to_unsigned(16#8A#, 8);
  gmul3_5(143) <= to_unsigned(16#AB#, 8);
  gmul3_5(144) <= to_unsigned(16#A8#, 8);
  gmul3_5(145) <= to_unsigned(16#AD#, 8);
  gmul3_5(146) <= to_unsigned(16#AE#, 8);
  gmul3_5(147) <= to_unsigned(16#A7#, 8);
  gmul3_5(148) <= to_unsigned(16#A4#, 8);
  gmul3_5(149) <= to_unsigned(16#A1#, 8);
  gmul3_5(150) <= to_unsigned(16#A2#, 8);
  gmul3_5(151) <= to_unsigned(16#B3#, 8);
  gmul3_5(152) <= to_unsigned(16#B0#, 8);
  gmul3_5(153) <= to_unsigned(16#B5#, 8);
  gmul3_5(154) <= to_unsigned(16#B6#, 8);
  gmul3_5(155) <= to_unsigned(16#BF#, 8);
  gmul3_5(156) <= to_unsigned(16#BC#, 8);
  gmul3_5(157) <= to_unsigned(16#B9#, 8);
  gmul3_5(158) <= to_unsigned(16#BA#, 8);
  gmul3_5(159) <= to_unsigned(16#FB#, 8);
  gmul3_5(160) <= to_unsigned(16#F8#, 8);
  gmul3_5(161) <= to_unsigned(16#FD#, 8);
  gmul3_5(162) <= to_unsigned(16#FE#, 8);
  gmul3_5(163) <= to_unsigned(16#F7#, 8);
  gmul3_5(164) <= to_unsigned(16#F4#, 8);
  gmul3_5(165) <= to_unsigned(16#F1#, 8);
  gmul3_5(166) <= to_unsigned(16#F2#, 8);
  gmul3_5(167) <= to_unsigned(16#E3#, 8);
  gmul3_5(168) <= to_unsigned(16#E0#, 8);
  gmul3_5(169) <= to_unsigned(16#E5#, 8);
  gmul3_5(170) <= to_unsigned(16#E6#, 8);
  gmul3_5(171) <= to_unsigned(16#EF#, 8);
  gmul3_5(172) <= to_unsigned(16#EC#, 8);
  gmul3_5(173) <= to_unsigned(16#E9#, 8);
  gmul3_5(174) <= to_unsigned(16#EA#, 8);
  gmul3_5(175) <= to_unsigned(16#CB#, 8);
  gmul3_5(176) <= to_unsigned(16#C8#, 8);
  gmul3_5(177) <= to_unsigned(16#CD#, 8);
  gmul3_5(178) <= to_unsigned(16#CE#, 8);
  gmul3_5(179) <= to_unsigned(16#C7#, 8);
  gmul3_5(180) <= to_unsigned(16#C4#, 8);
  gmul3_5(181) <= to_unsigned(16#C1#, 8);
  gmul3_5(182) <= to_unsigned(16#C2#, 8);
  gmul3_5(183) <= to_unsigned(16#D3#, 8);
  gmul3_5(184) <= to_unsigned(16#D0#, 8);
  gmul3_5(185) <= to_unsigned(16#D5#, 8);
  gmul3_5(186) <= to_unsigned(16#D6#, 8);
  gmul3_5(187) <= to_unsigned(16#DF#, 8);
  gmul3_5(188) <= to_unsigned(16#DC#, 8);
  gmul3_5(189) <= to_unsigned(16#D9#, 8);
  gmul3_5(190) <= to_unsigned(16#DA#, 8);
  gmul3_5(191) <= to_unsigned(16#5B#, 8);
  gmul3_5(192) <= to_unsigned(16#58#, 8);
  gmul3_5(193) <= to_unsigned(16#5D#, 8);
  gmul3_5(194) <= to_unsigned(16#5E#, 8);
  gmul3_5(195) <= to_unsigned(16#57#, 8);
  gmul3_5(196) <= to_unsigned(16#54#, 8);
  gmul3_5(197) <= to_unsigned(16#51#, 8);
  gmul3_5(198) <= to_unsigned(16#52#, 8);
  gmul3_5(199) <= to_unsigned(16#43#, 8);
  gmul3_5(200) <= to_unsigned(16#40#, 8);
  gmul3_5(201) <= to_unsigned(16#45#, 8);
  gmul3_5(202) <= to_unsigned(16#46#, 8);
  gmul3_5(203) <= to_unsigned(16#4F#, 8);
  gmul3_5(204) <= to_unsigned(16#4C#, 8);
  gmul3_5(205) <= to_unsigned(16#49#, 8);
  gmul3_5(206) <= to_unsigned(16#4A#, 8);
  gmul3_5(207) <= to_unsigned(16#6B#, 8);
  gmul3_5(208) <= to_unsigned(16#68#, 8);
  gmul3_5(209) <= to_unsigned(16#6D#, 8);
  gmul3_5(210) <= to_unsigned(16#6E#, 8);
  gmul3_5(211) <= to_unsigned(16#67#, 8);
  gmul3_5(212) <= to_unsigned(16#64#, 8);
  gmul3_5(213) <= to_unsigned(16#61#, 8);
  gmul3_5(214) <= to_unsigned(16#62#, 8);
  gmul3_5(215) <= to_unsigned(16#73#, 8);
  gmul3_5(216) <= to_unsigned(16#70#, 8);
  gmul3_5(217) <= to_unsigned(16#75#, 8);
  gmul3_5(218) <= to_unsigned(16#76#, 8);
  gmul3_5(219) <= to_unsigned(16#7F#, 8);
  gmul3_5(220) <= to_unsigned(16#7C#, 8);
  gmul3_5(221) <= to_unsigned(16#79#, 8);
  gmul3_5(222) <= to_unsigned(16#7A#, 8);
  gmul3_5(223) <= to_unsigned(16#3B#, 8);
  gmul3_5(224) <= to_unsigned(16#38#, 8);
  gmul3_5(225) <= to_unsigned(16#3D#, 8);
  gmul3_5(226) <= to_unsigned(16#3E#, 8);
  gmul3_5(227) <= to_unsigned(16#37#, 8);
  gmul3_5(228) <= to_unsigned(16#34#, 8);
  gmul3_5(229) <= to_unsigned(16#31#, 8);
  gmul3_5(230) <= to_unsigned(16#32#, 8);
  gmul3_5(231) <= to_unsigned(16#23#, 8);
  gmul3_5(232) <= to_unsigned(16#20#, 8);
  gmul3_5(233) <= to_unsigned(16#25#, 8);
  gmul3_5(234) <= to_unsigned(16#26#, 8);
  gmul3_5(235) <= to_unsigned(16#2F#, 8);
  gmul3_5(236) <= to_unsigned(16#2C#, 8);
  gmul3_5(237) <= to_unsigned(16#29#, 8);
  gmul3_5(238) <= to_unsigned(16#2A#, 8);
  gmul3_5(239) <= to_unsigned(16#0B#, 8);
  gmul3_5(240) <= to_unsigned(16#08#, 8);
  gmul3_5(241) <= to_unsigned(16#0D#, 8);
  gmul3_5(242) <= to_unsigned(16#0E#, 8);
  gmul3_5(243) <= to_unsigned(16#07#, 8);
  gmul3_5(244) <= to_unsigned(16#04#, 8);
  gmul3_5(245) <= to_unsigned(16#01#, 8);
  gmul3_5(246) <= to_unsigned(16#02#, 8);
  gmul3_5(247) <= to_unsigned(16#13#, 8);
  gmul3_5(248) <= to_unsigned(16#10#, 8);
  gmul3_5(249) <= to_unsigned(16#15#, 8);
  gmul3_5(250) <= to_unsigned(16#16#, 8);
  gmul3_5(251) <= to_unsigned(16#1F#, 8);
  gmul3_5(252) <= to_unsigned(16#1C#, 8);
  gmul3_5(253) <= to_unsigned(16#19#, 8);
  gmul3_5(254) <= to_unsigned(16#1A#, 8);
  gmul3_5(255) <= to_unsigned(16#1A#, 8);

  gmul2_6(0) <= to_unsigned(16#02#, 8);
  gmul2_6(1) <= to_unsigned(16#04#, 8);
  gmul2_6(2) <= to_unsigned(16#06#, 8);
  gmul2_6(3) <= to_unsigned(16#08#, 8);
  gmul2_6(4) <= to_unsigned(16#0A#, 8);
  gmul2_6(5) <= to_unsigned(16#0C#, 8);
  gmul2_6(6) <= to_unsigned(16#0E#, 8);
  gmul2_6(7) <= to_unsigned(16#10#, 8);
  gmul2_6(8) <= to_unsigned(16#12#, 8);
  gmul2_6(9) <= to_unsigned(16#14#, 8);
  gmul2_6(10) <= to_unsigned(16#16#, 8);
  gmul2_6(11) <= to_unsigned(16#18#, 8);
  gmul2_6(12) <= to_unsigned(16#1A#, 8);
  gmul2_6(13) <= to_unsigned(16#1C#, 8);
  gmul2_6(14) <= to_unsigned(16#1E#, 8);
  gmul2_6(15) <= to_unsigned(16#20#, 8);
  gmul2_6(16) <= to_unsigned(16#22#, 8);
  gmul2_6(17) <= to_unsigned(16#24#, 8);
  gmul2_6(18) <= to_unsigned(16#26#, 8);
  gmul2_6(19) <= to_unsigned(16#28#, 8);
  gmul2_6(20) <= to_unsigned(16#2A#, 8);
  gmul2_6(21) <= to_unsigned(16#2C#, 8);
  gmul2_6(22) <= to_unsigned(16#2E#, 8);
  gmul2_6(23) <= to_unsigned(16#30#, 8);
  gmul2_6(24) <= to_unsigned(16#32#, 8);
  gmul2_6(25) <= to_unsigned(16#34#, 8);
  gmul2_6(26) <= to_unsigned(16#36#, 8);
  gmul2_6(27) <= to_unsigned(16#38#, 8);
  gmul2_6(28) <= to_unsigned(16#3A#, 8);
  gmul2_6(29) <= to_unsigned(16#3C#, 8);
  gmul2_6(30) <= to_unsigned(16#3E#, 8);
  gmul2_6(31) <= to_unsigned(16#40#, 8);
  gmul2_6(32) <= to_unsigned(16#42#, 8);
  gmul2_6(33) <= to_unsigned(16#44#, 8);
  gmul2_6(34) <= to_unsigned(16#46#, 8);
  gmul2_6(35) <= to_unsigned(16#48#, 8);
  gmul2_6(36) <= to_unsigned(16#4A#, 8);
  gmul2_6(37) <= to_unsigned(16#4C#, 8);
  gmul2_6(38) <= to_unsigned(16#4E#, 8);
  gmul2_6(39) <= to_unsigned(16#50#, 8);
  gmul2_6(40) <= to_unsigned(16#52#, 8);
  gmul2_6(41) <= to_unsigned(16#54#, 8);
  gmul2_6(42) <= to_unsigned(16#56#, 8);
  gmul2_6(43) <= to_unsigned(16#58#, 8);
  gmul2_6(44) <= to_unsigned(16#5A#, 8);
  gmul2_6(45) <= to_unsigned(16#5C#, 8);
  gmul2_6(46) <= to_unsigned(16#5E#, 8);
  gmul2_6(47) <= to_unsigned(16#60#, 8);
  gmul2_6(48) <= to_unsigned(16#62#, 8);
  gmul2_6(49) <= to_unsigned(16#64#, 8);
  gmul2_6(50) <= to_unsigned(16#66#, 8);
  gmul2_6(51) <= to_unsigned(16#68#, 8);
  gmul2_6(52) <= to_unsigned(16#6A#, 8);
  gmul2_6(53) <= to_unsigned(16#6C#, 8);
  gmul2_6(54) <= to_unsigned(16#6E#, 8);
  gmul2_6(55) <= to_unsigned(16#70#, 8);
  gmul2_6(56) <= to_unsigned(16#72#, 8);
  gmul2_6(57) <= to_unsigned(16#74#, 8);
  gmul2_6(58) <= to_unsigned(16#76#, 8);
  gmul2_6(59) <= to_unsigned(16#78#, 8);
  gmul2_6(60) <= to_unsigned(16#7A#, 8);
  gmul2_6(61) <= to_unsigned(16#7C#, 8);
  gmul2_6(62) <= to_unsigned(16#7E#, 8);
  gmul2_6(63) <= to_unsigned(16#80#, 8);
  gmul2_6(64) <= to_unsigned(16#82#, 8);
  gmul2_6(65) <= to_unsigned(16#84#, 8);
  gmul2_6(66) <= to_unsigned(16#86#, 8);
  gmul2_6(67) <= to_unsigned(16#88#, 8);
  gmul2_6(68) <= to_unsigned(16#8A#, 8);
  gmul2_6(69) <= to_unsigned(16#8C#, 8);
  gmul2_6(70) <= to_unsigned(16#8E#, 8);
  gmul2_6(71) <= to_unsigned(16#90#, 8);
  gmul2_6(72) <= to_unsigned(16#92#, 8);
  gmul2_6(73) <= to_unsigned(16#94#, 8);
  gmul2_6(74) <= to_unsigned(16#96#, 8);
  gmul2_6(75) <= to_unsigned(16#98#, 8);
  gmul2_6(76) <= to_unsigned(16#9A#, 8);
  gmul2_6(77) <= to_unsigned(16#9C#, 8);
  gmul2_6(78) <= to_unsigned(16#9E#, 8);
  gmul2_6(79) <= to_unsigned(16#A0#, 8);
  gmul2_6(80) <= to_unsigned(16#A2#, 8);
  gmul2_6(81) <= to_unsigned(16#A4#, 8);
  gmul2_6(82) <= to_unsigned(16#A6#, 8);
  gmul2_6(83) <= to_unsigned(16#A8#, 8);
  gmul2_6(84) <= to_unsigned(16#AA#, 8);
  gmul2_6(85) <= to_unsigned(16#AC#, 8);
  gmul2_6(86) <= to_unsigned(16#AE#, 8);
  gmul2_6(87) <= to_unsigned(16#B0#, 8);
  gmul2_6(88) <= to_unsigned(16#B2#, 8);
  gmul2_6(89) <= to_unsigned(16#B4#, 8);
  gmul2_6(90) <= to_unsigned(16#B6#, 8);
  gmul2_6(91) <= to_unsigned(16#B8#, 8);
  gmul2_6(92) <= to_unsigned(16#BA#, 8);
  gmul2_6(93) <= to_unsigned(16#BC#, 8);
  gmul2_6(94) <= to_unsigned(16#BE#, 8);
  gmul2_6(95) <= to_unsigned(16#C0#, 8);
  gmul2_6(96) <= to_unsigned(16#C2#, 8);
  gmul2_6(97) <= to_unsigned(16#C4#, 8);
  gmul2_6(98) <= to_unsigned(16#C6#, 8);
  gmul2_6(99) <= to_unsigned(16#C8#, 8);
  gmul2_6(100) <= to_unsigned(16#CA#, 8);
  gmul2_6(101) <= to_unsigned(16#CC#, 8);
  gmul2_6(102) <= to_unsigned(16#CE#, 8);
  gmul2_6(103) <= to_unsigned(16#D0#, 8);
  gmul2_6(104) <= to_unsigned(16#D2#, 8);
  gmul2_6(105) <= to_unsigned(16#D4#, 8);
  gmul2_6(106) <= to_unsigned(16#D6#, 8);
  gmul2_6(107) <= to_unsigned(16#D8#, 8);
  gmul2_6(108) <= to_unsigned(16#DA#, 8);
  gmul2_6(109) <= to_unsigned(16#DC#, 8);
  gmul2_6(110) <= to_unsigned(16#DE#, 8);
  gmul2_6(111) <= to_unsigned(16#E0#, 8);
  gmul2_6(112) <= to_unsigned(16#E2#, 8);
  gmul2_6(113) <= to_unsigned(16#E4#, 8);
  gmul2_6(114) <= to_unsigned(16#E6#, 8);
  gmul2_6(115) <= to_unsigned(16#E8#, 8);
  gmul2_6(116) <= to_unsigned(16#EA#, 8);
  gmul2_6(117) <= to_unsigned(16#EC#, 8);
  gmul2_6(118) <= to_unsigned(16#EE#, 8);
  gmul2_6(119) <= to_unsigned(16#F0#, 8);
  gmul2_6(120) <= to_unsigned(16#F2#, 8);
  gmul2_6(121) <= to_unsigned(16#F4#, 8);
  gmul2_6(122) <= to_unsigned(16#F6#, 8);
  gmul2_6(123) <= to_unsigned(16#F8#, 8);
  gmul2_6(124) <= to_unsigned(16#FA#, 8);
  gmul2_6(125) <= to_unsigned(16#FC#, 8);
  gmul2_6(126) <= to_unsigned(16#FE#, 8);
  gmul2_6(127) <= to_unsigned(16#1B#, 8);
  gmul2_6(128) <= to_unsigned(16#19#, 8);
  gmul2_6(129) <= to_unsigned(16#1F#, 8);
  gmul2_6(130) <= to_unsigned(16#1D#, 8);
  gmul2_6(131) <= to_unsigned(16#13#, 8);
  gmul2_6(132) <= to_unsigned(16#11#, 8);
  gmul2_6(133) <= to_unsigned(16#17#, 8);
  gmul2_6(134) <= to_unsigned(16#15#, 8);
  gmul2_6(135) <= to_unsigned(16#0B#, 8);
  gmul2_6(136) <= to_unsigned(16#09#, 8);
  gmul2_6(137) <= to_unsigned(16#0F#, 8);
  gmul2_6(138) <= to_unsigned(16#0D#, 8);
  gmul2_6(139) <= to_unsigned(16#03#, 8);
  gmul2_6(140) <= to_unsigned(16#01#, 8);
  gmul2_6(141) <= to_unsigned(16#07#, 8);
  gmul2_6(142) <= to_unsigned(16#05#, 8);
  gmul2_6(143) <= to_unsigned(16#3B#, 8);
  gmul2_6(144) <= to_unsigned(16#39#, 8);
  gmul2_6(145) <= to_unsigned(16#3F#, 8);
  gmul2_6(146) <= to_unsigned(16#3D#, 8);
  gmul2_6(147) <= to_unsigned(16#33#, 8);
  gmul2_6(148) <= to_unsigned(16#31#, 8);
  gmul2_6(149) <= to_unsigned(16#37#, 8);
  gmul2_6(150) <= to_unsigned(16#35#, 8);
  gmul2_6(151) <= to_unsigned(16#2B#, 8);
  gmul2_6(152) <= to_unsigned(16#29#, 8);
  gmul2_6(153) <= to_unsigned(16#2F#, 8);
  gmul2_6(154) <= to_unsigned(16#2D#, 8);
  gmul2_6(155) <= to_unsigned(16#23#, 8);
  gmul2_6(156) <= to_unsigned(16#21#, 8);
  gmul2_6(157) <= to_unsigned(16#27#, 8);
  gmul2_6(158) <= to_unsigned(16#25#, 8);
  gmul2_6(159) <= to_unsigned(16#5B#, 8);
  gmul2_6(160) <= to_unsigned(16#59#, 8);
  gmul2_6(161) <= to_unsigned(16#5F#, 8);
  gmul2_6(162) <= to_unsigned(16#5D#, 8);
  gmul2_6(163) <= to_unsigned(16#53#, 8);
  gmul2_6(164) <= to_unsigned(16#51#, 8);
  gmul2_6(165) <= to_unsigned(16#57#, 8);
  gmul2_6(166) <= to_unsigned(16#55#, 8);
  gmul2_6(167) <= to_unsigned(16#4B#, 8);
  gmul2_6(168) <= to_unsigned(16#49#, 8);
  gmul2_6(169) <= to_unsigned(16#4F#, 8);
  gmul2_6(170) <= to_unsigned(16#4D#, 8);
  gmul2_6(171) <= to_unsigned(16#43#, 8);
  gmul2_6(172) <= to_unsigned(16#41#, 8);
  gmul2_6(173) <= to_unsigned(16#47#, 8);
  gmul2_6(174) <= to_unsigned(16#45#, 8);
  gmul2_6(175) <= to_unsigned(16#7B#, 8);
  gmul2_6(176) <= to_unsigned(16#79#, 8);
  gmul2_6(177) <= to_unsigned(16#7F#, 8);
  gmul2_6(178) <= to_unsigned(16#7D#, 8);
  gmul2_6(179) <= to_unsigned(16#73#, 8);
  gmul2_6(180) <= to_unsigned(16#71#, 8);
  gmul2_6(181) <= to_unsigned(16#77#, 8);
  gmul2_6(182) <= to_unsigned(16#75#, 8);
  gmul2_6(183) <= to_unsigned(16#6B#, 8);
  gmul2_6(184) <= to_unsigned(16#69#, 8);
  gmul2_6(185) <= to_unsigned(16#6F#, 8);
  gmul2_6(186) <= to_unsigned(16#6D#, 8);
  gmul2_6(187) <= to_unsigned(16#63#, 8);
  gmul2_6(188) <= to_unsigned(16#61#, 8);
  gmul2_6(189) <= to_unsigned(16#67#, 8);
  gmul2_6(190) <= to_unsigned(16#65#, 8);
  gmul2_6(191) <= to_unsigned(16#9B#, 8);
  gmul2_6(192) <= to_unsigned(16#99#, 8);
  gmul2_6(193) <= to_unsigned(16#9F#, 8);
  gmul2_6(194) <= to_unsigned(16#9D#, 8);
  gmul2_6(195) <= to_unsigned(16#93#, 8);
  gmul2_6(196) <= to_unsigned(16#91#, 8);
  gmul2_6(197) <= to_unsigned(16#97#, 8);
  gmul2_6(198) <= to_unsigned(16#95#, 8);
  gmul2_6(199) <= to_unsigned(16#8B#, 8);
  gmul2_6(200) <= to_unsigned(16#89#, 8);
  gmul2_6(201) <= to_unsigned(16#8F#, 8);
  gmul2_6(202) <= to_unsigned(16#8D#, 8);
  gmul2_6(203) <= to_unsigned(16#83#, 8);
  gmul2_6(204) <= to_unsigned(16#81#, 8);
  gmul2_6(205) <= to_unsigned(16#87#, 8);
  gmul2_6(206) <= to_unsigned(16#85#, 8);
  gmul2_6(207) <= to_unsigned(16#BB#, 8);
  gmul2_6(208) <= to_unsigned(16#B9#, 8);
  gmul2_6(209) <= to_unsigned(16#BF#, 8);
  gmul2_6(210) <= to_unsigned(16#BD#, 8);
  gmul2_6(211) <= to_unsigned(16#B3#, 8);
  gmul2_6(212) <= to_unsigned(16#B1#, 8);
  gmul2_6(213) <= to_unsigned(16#B7#, 8);
  gmul2_6(214) <= to_unsigned(16#B5#, 8);
  gmul2_6(215) <= to_unsigned(16#AB#, 8);
  gmul2_6(216) <= to_unsigned(16#A9#, 8);
  gmul2_6(217) <= to_unsigned(16#AF#, 8);
  gmul2_6(218) <= to_unsigned(16#AD#, 8);
  gmul2_6(219) <= to_unsigned(16#A3#, 8);
  gmul2_6(220) <= to_unsigned(16#A1#, 8);
  gmul2_6(221) <= to_unsigned(16#A7#, 8);
  gmul2_6(222) <= to_unsigned(16#A5#, 8);
  gmul2_6(223) <= to_unsigned(16#DB#, 8);
  gmul2_6(224) <= to_unsigned(16#D9#, 8);
  gmul2_6(225) <= to_unsigned(16#DF#, 8);
  gmul2_6(226) <= to_unsigned(16#DD#, 8);
  gmul2_6(227) <= to_unsigned(16#D3#, 8);
  gmul2_6(228) <= to_unsigned(16#D1#, 8);
  gmul2_6(229) <= to_unsigned(16#D7#, 8);
  gmul2_6(230) <= to_unsigned(16#D5#, 8);
  gmul2_6(231) <= to_unsigned(16#CB#, 8);
  gmul2_6(232) <= to_unsigned(16#C9#, 8);
  gmul2_6(233) <= to_unsigned(16#CF#, 8);
  gmul2_6(234) <= to_unsigned(16#CD#, 8);
  gmul2_6(235) <= to_unsigned(16#C3#, 8);
  gmul2_6(236) <= to_unsigned(16#C1#, 8);
  gmul2_6(237) <= to_unsigned(16#C7#, 8);
  gmul2_6(238) <= to_unsigned(16#C5#, 8);
  gmul2_6(239) <= to_unsigned(16#FB#, 8);
  gmul2_6(240) <= to_unsigned(16#F9#, 8);
  gmul2_6(241) <= to_unsigned(16#FF#, 8);
  gmul2_6(242) <= to_unsigned(16#FD#, 8);
  gmul2_6(243) <= to_unsigned(16#F3#, 8);
  gmul2_6(244) <= to_unsigned(16#F1#, 8);
  gmul2_6(245) <= to_unsigned(16#F7#, 8);
  gmul2_6(246) <= to_unsigned(16#F5#, 8);
  gmul2_6(247) <= to_unsigned(16#EB#, 8);
  gmul2_6(248) <= to_unsigned(16#E9#, 8);
  gmul2_6(249) <= to_unsigned(16#EF#, 8);
  gmul2_6(250) <= to_unsigned(16#ED#, 8);
  gmul2_6(251) <= to_unsigned(16#E3#, 8);
  gmul2_6(252) <= to_unsigned(16#E1#, 8);
  gmul2_6(253) <= to_unsigned(16#E7#, 8);
  gmul2_6(254) <= to_unsigned(16#E5#, 8);
  gmul2_6(255) <= to_unsigned(16#E5#, 8);

  gmul3_6(0) <= to_unsigned(16#03#, 8);
  gmul3_6(1) <= to_unsigned(16#06#, 8);
  gmul3_6(2) <= to_unsigned(16#05#, 8);
  gmul3_6(3) <= to_unsigned(16#0C#, 8);
  gmul3_6(4) <= to_unsigned(16#0F#, 8);
  gmul3_6(5) <= to_unsigned(16#0A#, 8);
  gmul3_6(6) <= to_unsigned(16#09#, 8);
  gmul3_6(7) <= to_unsigned(16#18#, 8);
  gmul3_6(8) <= to_unsigned(16#1B#, 8);
  gmul3_6(9) <= to_unsigned(16#1E#, 8);
  gmul3_6(10) <= to_unsigned(16#1D#, 8);
  gmul3_6(11) <= to_unsigned(16#14#, 8);
  gmul3_6(12) <= to_unsigned(16#17#, 8);
  gmul3_6(13) <= to_unsigned(16#12#, 8);
  gmul3_6(14) <= to_unsigned(16#11#, 8);
  gmul3_6(15) <= to_unsigned(16#30#, 8);
  gmul3_6(16) <= to_unsigned(16#33#, 8);
  gmul3_6(17) <= to_unsigned(16#36#, 8);
  gmul3_6(18) <= to_unsigned(16#35#, 8);
  gmul3_6(19) <= to_unsigned(16#3C#, 8);
  gmul3_6(20) <= to_unsigned(16#3F#, 8);
  gmul3_6(21) <= to_unsigned(16#3A#, 8);
  gmul3_6(22) <= to_unsigned(16#39#, 8);
  gmul3_6(23) <= to_unsigned(16#28#, 8);
  gmul3_6(24) <= to_unsigned(16#2B#, 8);
  gmul3_6(25) <= to_unsigned(16#2E#, 8);
  gmul3_6(26) <= to_unsigned(16#2D#, 8);
  gmul3_6(27) <= to_unsigned(16#24#, 8);
  gmul3_6(28) <= to_unsigned(16#27#, 8);
  gmul3_6(29) <= to_unsigned(16#22#, 8);
  gmul3_6(30) <= to_unsigned(16#21#, 8);
  gmul3_6(31) <= to_unsigned(16#60#, 8);
  gmul3_6(32) <= to_unsigned(16#63#, 8);
  gmul3_6(33) <= to_unsigned(16#66#, 8);
  gmul3_6(34) <= to_unsigned(16#65#, 8);
  gmul3_6(35) <= to_unsigned(16#6C#, 8);
  gmul3_6(36) <= to_unsigned(16#6F#, 8);
  gmul3_6(37) <= to_unsigned(16#6A#, 8);
  gmul3_6(38) <= to_unsigned(16#69#, 8);
  gmul3_6(39) <= to_unsigned(16#78#, 8);
  gmul3_6(40) <= to_unsigned(16#7B#, 8);
  gmul3_6(41) <= to_unsigned(16#7E#, 8);
  gmul3_6(42) <= to_unsigned(16#7D#, 8);
  gmul3_6(43) <= to_unsigned(16#74#, 8);
  gmul3_6(44) <= to_unsigned(16#77#, 8);
  gmul3_6(45) <= to_unsigned(16#72#, 8);
  gmul3_6(46) <= to_unsigned(16#71#, 8);
  gmul3_6(47) <= to_unsigned(16#50#, 8);
  gmul3_6(48) <= to_unsigned(16#53#, 8);
  gmul3_6(49) <= to_unsigned(16#56#, 8);
  gmul3_6(50) <= to_unsigned(16#55#, 8);
  gmul3_6(51) <= to_unsigned(16#5C#, 8);
  gmul3_6(52) <= to_unsigned(16#5F#, 8);
  gmul3_6(53) <= to_unsigned(16#5A#, 8);
  gmul3_6(54) <= to_unsigned(16#59#, 8);
  gmul3_6(55) <= to_unsigned(16#48#, 8);
  gmul3_6(56) <= to_unsigned(16#4B#, 8);
  gmul3_6(57) <= to_unsigned(16#4E#, 8);
  gmul3_6(58) <= to_unsigned(16#4D#, 8);
  gmul3_6(59) <= to_unsigned(16#44#, 8);
  gmul3_6(60) <= to_unsigned(16#47#, 8);
  gmul3_6(61) <= to_unsigned(16#42#, 8);
  gmul3_6(62) <= to_unsigned(16#41#, 8);
  gmul3_6(63) <= to_unsigned(16#C0#, 8);
  gmul3_6(64) <= to_unsigned(16#C3#, 8);
  gmul3_6(65) <= to_unsigned(16#C6#, 8);
  gmul3_6(66) <= to_unsigned(16#C5#, 8);
  gmul3_6(67) <= to_unsigned(16#CC#, 8);
  gmul3_6(68) <= to_unsigned(16#CF#, 8);
  gmul3_6(69) <= to_unsigned(16#CA#, 8);
  gmul3_6(70) <= to_unsigned(16#C9#, 8);
  gmul3_6(71) <= to_unsigned(16#D8#, 8);
  gmul3_6(72) <= to_unsigned(16#DB#, 8);
  gmul3_6(73) <= to_unsigned(16#DE#, 8);
  gmul3_6(74) <= to_unsigned(16#DD#, 8);
  gmul3_6(75) <= to_unsigned(16#D4#, 8);
  gmul3_6(76) <= to_unsigned(16#D7#, 8);
  gmul3_6(77) <= to_unsigned(16#D2#, 8);
  gmul3_6(78) <= to_unsigned(16#D1#, 8);
  gmul3_6(79) <= to_unsigned(16#F0#, 8);
  gmul3_6(80) <= to_unsigned(16#F3#, 8);
  gmul3_6(81) <= to_unsigned(16#F6#, 8);
  gmul3_6(82) <= to_unsigned(16#F5#, 8);
  gmul3_6(83) <= to_unsigned(16#FC#, 8);
  gmul3_6(84) <= to_unsigned(16#FF#, 8);
  gmul3_6(85) <= to_unsigned(16#FA#, 8);
  gmul3_6(86) <= to_unsigned(16#F9#, 8);
  gmul3_6(87) <= to_unsigned(16#E8#, 8);
  gmul3_6(88) <= to_unsigned(16#EB#, 8);
  gmul3_6(89) <= to_unsigned(16#EE#, 8);
  gmul3_6(90) <= to_unsigned(16#ED#, 8);
  gmul3_6(91) <= to_unsigned(16#E4#, 8);
  gmul3_6(92) <= to_unsigned(16#E7#, 8);
  gmul3_6(93) <= to_unsigned(16#E2#, 8);
  gmul3_6(94) <= to_unsigned(16#E1#, 8);
  gmul3_6(95) <= to_unsigned(16#A0#, 8);
  gmul3_6(96) <= to_unsigned(16#A3#, 8);
  gmul3_6(97) <= to_unsigned(16#A6#, 8);
  gmul3_6(98) <= to_unsigned(16#A5#, 8);
  gmul3_6(99) <= to_unsigned(16#AC#, 8);
  gmul3_6(100) <= to_unsigned(16#AF#, 8);
  gmul3_6(101) <= to_unsigned(16#AA#, 8);
  gmul3_6(102) <= to_unsigned(16#A9#, 8);
  gmul3_6(103) <= to_unsigned(16#B8#, 8);
  gmul3_6(104) <= to_unsigned(16#BB#, 8);
  gmul3_6(105) <= to_unsigned(16#BE#, 8);
  gmul3_6(106) <= to_unsigned(16#BD#, 8);
  gmul3_6(107) <= to_unsigned(16#B4#, 8);
  gmul3_6(108) <= to_unsigned(16#B7#, 8);
  gmul3_6(109) <= to_unsigned(16#B2#, 8);
  gmul3_6(110) <= to_unsigned(16#B1#, 8);
  gmul3_6(111) <= to_unsigned(16#90#, 8);
  gmul3_6(112) <= to_unsigned(16#93#, 8);
  gmul3_6(113) <= to_unsigned(16#96#, 8);
  gmul3_6(114) <= to_unsigned(16#95#, 8);
  gmul3_6(115) <= to_unsigned(16#9C#, 8);
  gmul3_6(116) <= to_unsigned(16#9F#, 8);
  gmul3_6(117) <= to_unsigned(16#9A#, 8);
  gmul3_6(118) <= to_unsigned(16#99#, 8);
  gmul3_6(119) <= to_unsigned(16#88#, 8);
  gmul3_6(120) <= to_unsigned(16#8B#, 8);
  gmul3_6(121) <= to_unsigned(16#8E#, 8);
  gmul3_6(122) <= to_unsigned(16#8D#, 8);
  gmul3_6(123) <= to_unsigned(16#84#, 8);
  gmul3_6(124) <= to_unsigned(16#87#, 8);
  gmul3_6(125) <= to_unsigned(16#82#, 8);
  gmul3_6(126) <= to_unsigned(16#81#, 8);
  gmul3_6(127) <= to_unsigned(16#9B#, 8);
  gmul3_6(128) <= to_unsigned(16#98#, 8);
  gmul3_6(129) <= to_unsigned(16#9D#, 8);
  gmul3_6(130) <= to_unsigned(16#9E#, 8);
  gmul3_6(131) <= to_unsigned(16#97#, 8);
  gmul3_6(132) <= to_unsigned(16#94#, 8);
  gmul3_6(133) <= to_unsigned(16#91#, 8);
  gmul3_6(134) <= to_unsigned(16#92#, 8);
  gmul3_6(135) <= to_unsigned(16#83#, 8);
  gmul3_6(136) <= to_unsigned(16#80#, 8);
  gmul3_6(137) <= to_unsigned(16#85#, 8);
  gmul3_6(138) <= to_unsigned(16#86#, 8);
  gmul3_6(139) <= to_unsigned(16#8F#, 8);
  gmul3_6(140) <= to_unsigned(16#8C#, 8);
  gmul3_6(141) <= to_unsigned(16#89#, 8);
  gmul3_6(142) <= to_unsigned(16#8A#, 8);
  gmul3_6(143) <= to_unsigned(16#AB#, 8);
  gmul3_6(144) <= to_unsigned(16#A8#, 8);
  gmul3_6(145) <= to_unsigned(16#AD#, 8);
  gmul3_6(146) <= to_unsigned(16#AE#, 8);
  gmul3_6(147) <= to_unsigned(16#A7#, 8);
  gmul3_6(148) <= to_unsigned(16#A4#, 8);
  gmul3_6(149) <= to_unsigned(16#A1#, 8);
  gmul3_6(150) <= to_unsigned(16#A2#, 8);
  gmul3_6(151) <= to_unsigned(16#B3#, 8);
  gmul3_6(152) <= to_unsigned(16#B0#, 8);
  gmul3_6(153) <= to_unsigned(16#B5#, 8);
  gmul3_6(154) <= to_unsigned(16#B6#, 8);
  gmul3_6(155) <= to_unsigned(16#BF#, 8);
  gmul3_6(156) <= to_unsigned(16#BC#, 8);
  gmul3_6(157) <= to_unsigned(16#B9#, 8);
  gmul3_6(158) <= to_unsigned(16#BA#, 8);
  gmul3_6(159) <= to_unsigned(16#FB#, 8);
  gmul3_6(160) <= to_unsigned(16#F8#, 8);
  gmul3_6(161) <= to_unsigned(16#FD#, 8);
  gmul3_6(162) <= to_unsigned(16#FE#, 8);
  gmul3_6(163) <= to_unsigned(16#F7#, 8);
  gmul3_6(164) <= to_unsigned(16#F4#, 8);
  gmul3_6(165) <= to_unsigned(16#F1#, 8);
  gmul3_6(166) <= to_unsigned(16#F2#, 8);
  gmul3_6(167) <= to_unsigned(16#E3#, 8);
  gmul3_6(168) <= to_unsigned(16#E0#, 8);
  gmul3_6(169) <= to_unsigned(16#E5#, 8);
  gmul3_6(170) <= to_unsigned(16#E6#, 8);
  gmul3_6(171) <= to_unsigned(16#EF#, 8);
  gmul3_6(172) <= to_unsigned(16#EC#, 8);
  gmul3_6(173) <= to_unsigned(16#E9#, 8);
  gmul3_6(174) <= to_unsigned(16#EA#, 8);
  gmul3_6(175) <= to_unsigned(16#CB#, 8);
  gmul3_6(176) <= to_unsigned(16#C8#, 8);
  gmul3_6(177) <= to_unsigned(16#CD#, 8);
  gmul3_6(178) <= to_unsigned(16#CE#, 8);
  gmul3_6(179) <= to_unsigned(16#C7#, 8);
  gmul3_6(180) <= to_unsigned(16#C4#, 8);
  gmul3_6(181) <= to_unsigned(16#C1#, 8);
  gmul3_6(182) <= to_unsigned(16#C2#, 8);
  gmul3_6(183) <= to_unsigned(16#D3#, 8);
  gmul3_6(184) <= to_unsigned(16#D0#, 8);
  gmul3_6(185) <= to_unsigned(16#D5#, 8);
  gmul3_6(186) <= to_unsigned(16#D6#, 8);
  gmul3_6(187) <= to_unsigned(16#DF#, 8);
  gmul3_6(188) <= to_unsigned(16#DC#, 8);
  gmul3_6(189) <= to_unsigned(16#D9#, 8);
  gmul3_6(190) <= to_unsigned(16#DA#, 8);
  gmul3_6(191) <= to_unsigned(16#5B#, 8);
  gmul3_6(192) <= to_unsigned(16#58#, 8);
  gmul3_6(193) <= to_unsigned(16#5D#, 8);
  gmul3_6(194) <= to_unsigned(16#5E#, 8);
  gmul3_6(195) <= to_unsigned(16#57#, 8);
  gmul3_6(196) <= to_unsigned(16#54#, 8);
  gmul3_6(197) <= to_unsigned(16#51#, 8);
  gmul3_6(198) <= to_unsigned(16#52#, 8);
  gmul3_6(199) <= to_unsigned(16#43#, 8);
  gmul3_6(200) <= to_unsigned(16#40#, 8);
  gmul3_6(201) <= to_unsigned(16#45#, 8);
  gmul3_6(202) <= to_unsigned(16#46#, 8);
  gmul3_6(203) <= to_unsigned(16#4F#, 8);
  gmul3_6(204) <= to_unsigned(16#4C#, 8);
  gmul3_6(205) <= to_unsigned(16#49#, 8);
  gmul3_6(206) <= to_unsigned(16#4A#, 8);
  gmul3_6(207) <= to_unsigned(16#6B#, 8);
  gmul3_6(208) <= to_unsigned(16#68#, 8);
  gmul3_6(209) <= to_unsigned(16#6D#, 8);
  gmul3_6(210) <= to_unsigned(16#6E#, 8);
  gmul3_6(211) <= to_unsigned(16#67#, 8);
  gmul3_6(212) <= to_unsigned(16#64#, 8);
  gmul3_6(213) <= to_unsigned(16#61#, 8);
  gmul3_6(214) <= to_unsigned(16#62#, 8);
  gmul3_6(215) <= to_unsigned(16#73#, 8);
  gmul3_6(216) <= to_unsigned(16#70#, 8);
  gmul3_6(217) <= to_unsigned(16#75#, 8);
  gmul3_6(218) <= to_unsigned(16#76#, 8);
  gmul3_6(219) <= to_unsigned(16#7F#, 8);
  gmul3_6(220) <= to_unsigned(16#7C#, 8);
  gmul3_6(221) <= to_unsigned(16#79#, 8);
  gmul3_6(222) <= to_unsigned(16#7A#, 8);
  gmul3_6(223) <= to_unsigned(16#3B#, 8);
  gmul3_6(224) <= to_unsigned(16#38#, 8);
  gmul3_6(225) <= to_unsigned(16#3D#, 8);
  gmul3_6(226) <= to_unsigned(16#3E#, 8);
  gmul3_6(227) <= to_unsigned(16#37#, 8);
  gmul3_6(228) <= to_unsigned(16#34#, 8);
  gmul3_6(229) <= to_unsigned(16#31#, 8);
  gmul3_6(230) <= to_unsigned(16#32#, 8);
  gmul3_6(231) <= to_unsigned(16#23#, 8);
  gmul3_6(232) <= to_unsigned(16#20#, 8);
  gmul3_6(233) <= to_unsigned(16#25#, 8);
  gmul3_6(234) <= to_unsigned(16#26#, 8);
  gmul3_6(235) <= to_unsigned(16#2F#, 8);
  gmul3_6(236) <= to_unsigned(16#2C#, 8);
  gmul3_6(237) <= to_unsigned(16#29#, 8);
  gmul3_6(238) <= to_unsigned(16#2A#, 8);
  gmul3_6(239) <= to_unsigned(16#0B#, 8);
  gmul3_6(240) <= to_unsigned(16#08#, 8);
  gmul3_6(241) <= to_unsigned(16#0D#, 8);
  gmul3_6(242) <= to_unsigned(16#0E#, 8);
  gmul3_6(243) <= to_unsigned(16#07#, 8);
  gmul3_6(244) <= to_unsigned(16#04#, 8);
  gmul3_6(245) <= to_unsigned(16#01#, 8);
  gmul3_6(246) <= to_unsigned(16#02#, 8);
  gmul3_6(247) <= to_unsigned(16#13#, 8);
  gmul3_6(248) <= to_unsigned(16#10#, 8);
  gmul3_6(249) <= to_unsigned(16#15#, 8);
  gmul3_6(250) <= to_unsigned(16#16#, 8);
  gmul3_6(251) <= to_unsigned(16#1F#, 8);
  gmul3_6(252) <= to_unsigned(16#1C#, 8);
  gmul3_6(253) <= to_unsigned(16#19#, 8);
  gmul3_6(254) <= to_unsigned(16#1A#, 8);
  gmul3_6(255) <= to_unsigned(16#1A#, 8);

  gmul3_7(0) <= to_unsigned(16#03#, 8);
  gmul3_7(1) <= to_unsigned(16#06#, 8);
  gmul3_7(2) <= to_unsigned(16#05#, 8);
  gmul3_7(3) <= to_unsigned(16#0C#, 8);
  gmul3_7(4) <= to_unsigned(16#0F#, 8);
  gmul3_7(5) <= to_unsigned(16#0A#, 8);
  gmul3_7(6) <= to_unsigned(16#09#, 8);
  gmul3_7(7) <= to_unsigned(16#18#, 8);
  gmul3_7(8) <= to_unsigned(16#1B#, 8);
  gmul3_7(9) <= to_unsigned(16#1E#, 8);
  gmul3_7(10) <= to_unsigned(16#1D#, 8);
  gmul3_7(11) <= to_unsigned(16#14#, 8);
  gmul3_7(12) <= to_unsigned(16#17#, 8);
  gmul3_7(13) <= to_unsigned(16#12#, 8);
  gmul3_7(14) <= to_unsigned(16#11#, 8);
  gmul3_7(15) <= to_unsigned(16#30#, 8);
  gmul3_7(16) <= to_unsigned(16#33#, 8);
  gmul3_7(17) <= to_unsigned(16#36#, 8);
  gmul3_7(18) <= to_unsigned(16#35#, 8);
  gmul3_7(19) <= to_unsigned(16#3C#, 8);
  gmul3_7(20) <= to_unsigned(16#3F#, 8);
  gmul3_7(21) <= to_unsigned(16#3A#, 8);
  gmul3_7(22) <= to_unsigned(16#39#, 8);
  gmul3_7(23) <= to_unsigned(16#28#, 8);
  gmul3_7(24) <= to_unsigned(16#2B#, 8);
  gmul3_7(25) <= to_unsigned(16#2E#, 8);
  gmul3_7(26) <= to_unsigned(16#2D#, 8);
  gmul3_7(27) <= to_unsigned(16#24#, 8);
  gmul3_7(28) <= to_unsigned(16#27#, 8);
  gmul3_7(29) <= to_unsigned(16#22#, 8);
  gmul3_7(30) <= to_unsigned(16#21#, 8);
  gmul3_7(31) <= to_unsigned(16#60#, 8);
  gmul3_7(32) <= to_unsigned(16#63#, 8);
  gmul3_7(33) <= to_unsigned(16#66#, 8);
  gmul3_7(34) <= to_unsigned(16#65#, 8);
  gmul3_7(35) <= to_unsigned(16#6C#, 8);
  gmul3_7(36) <= to_unsigned(16#6F#, 8);
  gmul3_7(37) <= to_unsigned(16#6A#, 8);
  gmul3_7(38) <= to_unsigned(16#69#, 8);
  gmul3_7(39) <= to_unsigned(16#78#, 8);
  gmul3_7(40) <= to_unsigned(16#7B#, 8);
  gmul3_7(41) <= to_unsigned(16#7E#, 8);
  gmul3_7(42) <= to_unsigned(16#7D#, 8);
  gmul3_7(43) <= to_unsigned(16#74#, 8);
  gmul3_7(44) <= to_unsigned(16#77#, 8);
  gmul3_7(45) <= to_unsigned(16#72#, 8);
  gmul3_7(46) <= to_unsigned(16#71#, 8);
  gmul3_7(47) <= to_unsigned(16#50#, 8);
  gmul3_7(48) <= to_unsigned(16#53#, 8);
  gmul3_7(49) <= to_unsigned(16#56#, 8);
  gmul3_7(50) <= to_unsigned(16#55#, 8);
  gmul3_7(51) <= to_unsigned(16#5C#, 8);
  gmul3_7(52) <= to_unsigned(16#5F#, 8);
  gmul3_7(53) <= to_unsigned(16#5A#, 8);
  gmul3_7(54) <= to_unsigned(16#59#, 8);
  gmul3_7(55) <= to_unsigned(16#48#, 8);
  gmul3_7(56) <= to_unsigned(16#4B#, 8);
  gmul3_7(57) <= to_unsigned(16#4E#, 8);
  gmul3_7(58) <= to_unsigned(16#4D#, 8);
  gmul3_7(59) <= to_unsigned(16#44#, 8);
  gmul3_7(60) <= to_unsigned(16#47#, 8);
  gmul3_7(61) <= to_unsigned(16#42#, 8);
  gmul3_7(62) <= to_unsigned(16#41#, 8);
  gmul3_7(63) <= to_unsigned(16#C0#, 8);
  gmul3_7(64) <= to_unsigned(16#C3#, 8);
  gmul3_7(65) <= to_unsigned(16#C6#, 8);
  gmul3_7(66) <= to_unsigned(16#C5#, 8);
  gmul3_7(67) <= to_unsigned(16#CC#, 8);
  gmul3_7(68) <= to_unsigned(16#CF#, 8);
  gmul3_7(69) <= to_unsigned(16#CA#, 8);
  gmul3_7(70) <= to_unsigned(16#C9#, 8);
  gmul3_7(71) <= to_unsigned(16#D8#, 8);
  gmul3_7(72) <= to_unsigned(16#DB#, 8);
  gmul3_7(73) <= to_unsigned(16#DE#, 8);
  gmul3_7(74) <= to_unsigned(16#DD#, 8);
  gmul3_7(75) <= to_unsigned(16#D4#, 8);
  gmul3_7(76) <= to_unsigned(16#D7#, 8);
  gmul3_7(77) <= to_unsigned(16#D2#, 8);
  gmul3_7(78) <= to_unsigned(16#D1#, 8);
  gmul3_7(79) <= to_unsigned(16#F0#, 8);
  gmul3_7(80) <= to_unsigned(16#F3#, 8);
  gmul3_7(81) <= to_unsigned(16#F6#, 8);
  gmul3_7(82) <= to_unsigned(16#F5#, 8);
  gmul3_7(83) <= to_unsigned(16#FC#, 8);
  gmul3_7(84) <= to_unsigned(16#FF#, 8);
  gmul3_7(85) <= to_unsigned(16#FA#, 8);
  gmul3_7(86) <= to_unsigned(16#F9#, 8);
  gmul3_7(87) <= to_unsigned(16#E8#, 8);
  gmul3_7(88) <= to_unsigned(16#EB#, 8);
  gmul3_7(89) <= to_unsigned(16#EE#, 8);
  gmul3_7(90) <= to_unsigned(16#ED#, 8);
  gmul3_7(91) <= to_unsigned(16#E4#, 8);
  gmul3_7(92) <= to_unsigned(16#E7#, 8);
  gmul3_7(93) <= to_unsigned(16#E2#, 8);
  gmul3_7(94) <= to_unsigned(16#E1#, 8);
  gmul3_7(95) <= to_unsigned(16#A0#, 8);
  gmul3_7(96) <= to_unsigned(16#A3#, 8);
  gmul3_7(97) <= to_unsigned(16#A6#, 8);
  gmul3_7(98) <= to_unsigned(16#A5#, 8);
  gmul3_7(99) <= to_unsigned(16#AC#, 8);
  gmul3_7(100) <= to_unsigned(16#AF#, 8);
  gmul3_7(101) <= to_unsigned(16#AA#, 8);
  gmul3_7(102) <= to_unsigned(16#A9#, 8);
  gmul3_7(103) <= to_unsigned(16#B8#, 8);
  gmul3_7(104) <= to_unsigned(16#BB#, 8);
  gmul3_7(105) <= to_unsigned(16#BE#, 8);
  gmul3_7(106) <= to_unsigned(16#BD#, 8);
  gmul3_7(107) <= to_unsigned(16#B4#, 8);
  gmul3_7(108) <= to_unsigned(16#B7#, 8);
  gmul3_7(109) <= to_unsigned(16#B2#, 8);
  gmul3_7(110) <= to_unsigned(16#B1#, 8);
  gmul3_7(111) <= to_unsigned(16#90#, 8);
  gmul3_7(112) <= to_unsigned(16#93#, 8);
  gmul3_7(113) <= to_unsigned(16#96#, 8);
  gmul3_7(114) <= to_unsigned(16#95#, 8);
  gmul3_7(115) <= to_unsigned(16#9C#, 8);
  gmul3_7(116) <= to_unsigned(16#9F#, 8);
  gmul3_7(117) <= to_unsigned(16#9A#, 8);
  gmul3_7(118) <= to_unsigned(16#99#, 8);
  gmul3_7(119) <= to_unsigned(16#88#, 8);
  gmul3_7(120) <= to_unsigned(16#8B#, 8);
  gmul3_7(121) <= to_unsigned(16#8E#, 8);
  gmul3_7(122) <= to_unsigned(16#8D#, 8);
  gmul3_7(123) <= to_unsigned(16#84#, 8);
  gmul3_7(124) <= to_unsigned(16#87#, 8);
  gmul3_7(125) <= to_unsigned(16#82#, 8);
  gmul3_7(126) <= to_unsigned(16#81#, 8);
  gmul3_7(127) <= to_unsigned(16#9B#, 8);
  gmul3_7(128) <= to_unsigned(16#98#, 8);
  gmul3_7(129) <= to_unsigned(16#9D#, 8);
  gmul3_7(130) <= to_unsigned(16#9E#, 8);
  gmul3_7(131) <= to_unsigned(16#97#, 8);
  gmul3_7(132) <= to_unsigned(16#94#, 8);
  gmul3_7(133) <= to_unsigned(16#91#, 8);
  gmul3_7(134) <= to_unsigned(16#92#, 8);
  gmul3_7(135) <= to_unsigned(16#83#, 8);
  gmul3_7(136) <= to_unsigned(16#80#, 8);
  gmul3_7(137) <= to_unsigned(16#85#, 8);
  gmul3_7(138) <= to_unsigned(16#86#, 8);
  gmul3_7(139) <= to_unsigned(16#8F#, 8);
  gmul3_7(140) <= to_unsigned(16#8C#, 8);
  gmul3_7(141) <= to_unsigned(16#89#, 8);
  gmul3_7(142) <= to_unsigned(16#8A#, 8);
  gmul3_7(143) <= to_unsigned(16#AB#, 8);
  gmul3_7(144) <= to_unsigned(16#A8#, 8);
  gmul3_7(145) <= to_unsigned(16#AD#, 8);
  gmul3_7(146) <= to_unsigned(16#AE#, 8);
  gmul3_7(147) <= to_unsigned(16#A7#, 8);
  gmul3_7(148) <= to_unsigned(16#A4#, 8);
  gmul3_7(149) <= to_unsigned(16#A1#, 8);
  gmul3_7(150) <= to_unsigned(16#A2#, 8);
  gmul3_7(151) <= to_unsigned(16#B3#, 8);
  gmul3_7(152) <= to_unsigned(16#B0#, 8);
  gmul3_7(153) <= to_unsigned(16#B5#, 8);
  gmul3_7(154) <= to_unsigned(16#B6#, 8);
  gmul3_7(155) <= to_unsigned(16#BF#, 8);
  gmul3_7(156) <= to_unsigned(16#BC#, 8);
  gmul3_7(157) <= to_unsigned(16#B9#, 8);
  gmul3_7(158) <= to_unsigned(16#BA#, 8);
  gmul3_7(159) <= to_unsigned(16#FB#, 8);
  gmul3_7(160) <= to_unsigned(16#F8#, 8);
  gmul3_7(161) <= to_unsigned(16#FD#, 8);
  gmul3_7(162) <= to_unsigned(16#FE#, 8);
  gmul3_7(163) <= to_unsigned(16#F7#, 8);
  gmul3_7(164) <= to_unsigned(16#F4#, 8);
  gmul3_7(165) <= to_unsigned(16#F1#, 8);
  gmul3_7(166) <= to_unsigned(16#F2#, 8);
  gmul3_7(167) <= to_unsigned(16#E3#, 8);
  gmul3_7(168) <= to_unsigned(16#E0#, 8);
  gmul3_7(169) <= to_unsigned(16#E5#, 8);
  gmul3_7(170) <= to_unsigned(16#E6#, 8);
  gmul3_7(171) <= to_unsigned(16#EF#, 8);
  gmul3_7(172) <= to_unsigned(16#EC#, 8);
  gmul3_7(173) <= to_unsigned(16#E9#, 8);
  gmul3_7(174) <= to_unsigned(16#EA#, 8);
  gmul3_7(175) <= to_unsigned(16#CB#, 8);
  gmul3_7(176) <= to_unsigned(16#C8#, 8);
  gmul3_7(177) <= to_unsigned(16#CD#, 8);
  gmul3_7(178) <= to_unsigned(16#CE#, 8);
  gmul3_7(179) <= to_unsigned(16#C7#, 8);
  gmul3_7(180) <= to_unsigned(16#C4#, 8);
  gmul3_7(181) <= to_unsigned(16#C1#, 8);
  gmul3_7(182) <= to_unsigned(16#C2#, 8);
  gmul3_7(183) <= to_unsigned(16#D3#, 8);
  gmul3_7(184) <= to_unsigned(16#D0#, 8);
  gmul3_7(185) <= to_unsigned(16#D5#, 8);
  gmul3_7(186) <= to_unsigned(16#D6#, 8);
  gmul3_7(187) <= to_unsigned(16#DF#, 8);
  gmul3_7(188) <= to_unsigned(16#DC#, 8);
  gmul3_7(189) <= to_unsigned(16#D9#, 8);
  gmul3_7(190) <= to_unsigned(16#DA#, 8);
  gmul3_7(191) <= to_unsigned(16#5B#, 8);
  gmul3_7(192) <= to_unsigned(16#58#, 8);
  gmul3_7(193) <= to_unsigned(16#5D#, 8);
  gmul3_7(194) <= to_unsigned(16#5E#, 8);
  gmul3_7(195) <= to_unsigned(16#57#, 8);
  gmul3_7(196) <= to_unsigned(16#54#, 8);
  gmul3_7(197) <= to_unsigned(16#51#, 8);
  gmul3_7(198) <= to_unsigned(16#52#, 8);
  gmul3_7(199) <= to_unsigned(16#43#, 8);
  gmul3_7(200) <= to_unsigned(16#40#, 8);
  gmul3_7(201) <= to_unsigned(16#45#, 8);
  gmul3_7(202) <= to_unsigned(16#46#, 8);
  gmul3_7(203) <= to_unsigned(16#4F#, 8);
  gmul3_7(204) <= to_unsigned(16#4C#, 8);
  gmul3_7(205) <= to_unsigned(16#49#, 8);
  gmul3_7(206) <= to_unsigned(16#4A#, 8);
  gmul3_7(207) <= to_unsigned(16#6B#, 8);
  gmul3_7(208) <= to_unsigned(16#68#, 8);
  gmul3_7(209) <= to_unsigned(16#6D#, 8);
  gmul3_7(210) <= to_unsigned(16#6E#, 8);
  gmul3_7(211) <= to_unsigned(16#67#, 8);
  gmul3_7(212) <= to_unsigned(16#64#, 8);
  gmul3_7(213) <= to_unsigned(16#61#, 8);
  gmul3_7(214) <= to_unsigned(16#62#, 8);
  gmul3_7(215) <= to_unsigned(16#73#, 8);
  gmul3_7(216) <= to_unsigned(16#70#, 8);
  gmul3_7(217) <= to_unsigned(16#75#, 8);
  gmul3_7(218) <= to_unsigned(16#76#, 8);
  gmul3_7(219) <= to_unsigned(16#7F#, 8);
  gmul3_7(220) <= to_unsigned(16#7C#, 8);
  gmul3_7(221) <= to_unsigned(16#79#, 8);
  gmul3_7(222) <= to_unsigned(16#7A#, 8);
  gmul3_7(223) <= to_unsigned(16#3B#, 8);
  gmul3_7(224) <= to_unsigned(16#38#, 8);
  gmul3_7(225) <= to_unsigned(16#3D#, 8);
  gmul3_7(226) <= to_unsigned(16#3E#, 8);
  gmul3_7(227) <= to_unsigned(16#37#, 8);
  gmul3_7(228) <= to_unsigned(16#34#, 8);
  gmul3_7(229) <= to_unsigned(16#31#, 8);
  gmul3_7(230) <= to_unsigned(16#32#, 8);
  gmul3_7(231) <= to_unsigned(16#23#, 8);
  gmul3_7(232) <= to_unsigned(16#20#, 8);
  gmul3_7(233) <= to_unsigned(16#25#, 8);
  gmul3_7(234) <= to_unsigned(16#26#, 8);
  gmul3_7(235) <= to_unsigned(16#2F#, 8);
  gmul3_7(236) <= to_unsigned(16#2C#, 8);
  gmul3_7(237) <= to_unsigned(16#29#, 8);
  gmul3_7(238) <= to_unsigned(16#2A#, 8);
  gmul3_7(239) <= to_unsigned(16#0B#, 8);
  gmul3_7(240) <= to_unsigned(16#08#, 8);
  gmul3_7(241) <= to_unsigned(16#0D#, 8);
  gmul3_7(242) <= to_unsigned(16#0E#, 8);
  gmul3_7(243) <= to_unsigned(16#07#, 8);
  gmul3_7(244) <= to_unsigned(16#04#, 8);
  gmul3_7(245) <= to_unsigned(16#01#, 8);
  gmul3_7(246) <= to_unsigned(16#02#, 8);
  gmul3_7(247) <= to_unsigned(16#13#, 8);
  gmul3_7(248) <= to_unsigned(16#10#, 8);
  gmul3_7(249) <= to_unsigned(16#15#, 8);
  gmul3_7(250) <= to_unsigned(16#16#, 8);
  gmul3_7(251) <= to_unsigned(16#1F#, 8);
  gmul3_7(252) <= to_unsigned(16#1C#, 8);
  gmul3_7(253) <= to_unsigned(16#19#, 8);
  gmul3_7(254) <= to_unsigned(16#1A#, 8);
  gmul3_7(255) <= to_unsigned(16#1A#, 8);

  gmul2_7(0) <= to_unsigned(16#02#, 8);
  gmul2_7(1) <= to_unsigned(16#04#, 8);
  gmul2_7(2) <= to_unsigned(16#06#, 8);
  gmul2_7(3) <= to_unsigned(16#08#, 8);
  gmul2_7(4) <= to_unsigned(16#0A#, 8);
  gmul2_7(5) <= to_unsigned(16#0C#, 8);
  gmul2_7(6) <= to_unsigned(16#0E#, 8);
  gmul2_7(7) <= to_unsigned(16#10#, 8);
  gmul2_7(8) <= to_unsigned(16#12#, 8);
  gmul2_7(9) <= to_unsigned(16#14#, 8);
  gmul2_7(10) <= to_unsigned(16#16#, 8);
  gmul2_7(11) <= to_unsigned(16#18#, 8);
  gmul2_7(12) <= to_unsigned(16#1A#, 8);
  gmul2_7(13) <= to_unsigned(16#1C#, 8);
  gmul2_7(14) <= to_unsigned(16#1E#, 8);
  gmul2_7(15) <= to_unsigned(16#20#, 8);
  gmul2_7(16) <= to_unsigned(16#22#, 8);
  gmul2_7(17) <= to_unsigned(16#24#, 8);
  gmul2_7(18) <= to_unsigned(16#26#, 8);
  gmul2_7(19) <= to_unsigned(16#28#, 8);
  gmul2_7(20) <= to_unsigned(16#2A#, 8);
  gmul2_7(21) <= to_unsigned(16#2C#, 8);
  gmul2_7(22) <= to_unsigned(16#2E#, 8);
  gmul2_7(23) <= to_unsigned(16#30#, 8);
  gmul2_7(24) <= to_unsigned(16#32#, 8);
  gmul2_7(25) <= to_unsigned(16#34#, 8);
  gmul2_7(26) <= to_unsigned(16#36#, 8);
  gmul2_7(27) <= to_unsigned(16#38#, 8);
  gmul2_7(28) <= to_unsigned(16#3A#, 8);
  gmul2_7(29) <= to_unsigned(16#3C#, 8);
  gmul2_7(30) <= to_unsigned(16#3E#, 8);
  gmul2_7(31) <= to_unsigned(16#40#, 8);
  gmul2_7(32) <= to_unsigned(16#42#, 8);
  gmul2_7(33) <= to_unsigned(16#44#, 8);
  gmul2_7(34) <= to_unsigned(16#46#, 8);
  gmul2_7(35) <= to_unsigned(16#48#, 8);
  gmul2_7(36) <= to_unsigned(16#4A#, 8);
  gmul2_7(37) <= to_unsigned(16#4C#, 8);
  gmul2_7(38) <= to_unsigned(16#4E#, 8);
  gmul2_7(39) <= to_unsigned(16#50#, 8);
  gmul2_7(40) <= to_unsigned(16#52#, 8);
  gmul2_7(41) <= to_unsigned(16#54#, 8);
  gmul2_7(42) <= to_unsigned(16#56#, 8);
  gmul2_7(43) <= to_unsigned(16#58#, 8);
  gmul2_7(44) <= to_unsigned(16#5A#, 8);
  gmul2_7(45) <= to_unsigned(16#5C#, 8);
  gmul2_7(46) <= to_unsigned(16#5E#, 8);
  gmul2_7(47) <= to_unsigned(16#60#, 8);
  gmul2_7(48) <= to_unsigned(16#62#, 8);
  gmul2_7(49) <= to_unsigned(16#64#, 8);
  gmul2_7(50) <= to_unsigned(16#66#, 8);
  gmul2_7(51) <= to_unsigned(16#68#, 8);
  gmul2_7(52) <= to_unsigned(16#6A#, 8);
  gmul2_7(53) <= to_unsigned(16#6C#, 8);
  gmul2_7(54) <= to_unsigned(16#6E#, 8);
  gmul2_7(55) <= to_unsigned(16#70#, 8);
  gmul2_7(56) <= to_unsigned(16#72#, 8);
  gmul2_7(57) <= to_unsigned(16#74#, 8);
  gmul2_7(58) <= to_unsigned(16#76#, 8);
  gmul2_7(59) <= to_unsigned(16#78#, 8);
  gmul2_7(60) <= to_unsigned(16#7A#, 8);
  gmul2_7(61) <= to_unsigned(16#7C#, 8);
  gmul2_7(62) <= to_unsigned(16#7E#, 8);
  gmul2_7(63) <= to_unsigned(16#80#, 8);
  gmul2_7(64) <= to_unsigned(16#82#, 8);
  gmul2_7(65) <= to_unsigned(16#84#, 8);
  gmul2_7(66) <= to_unsigned(16#86#, 8);
  gmul2_7(67) <= to_unsigned(16#88#, 8);
  gmul2_7(68) <= to_unsigned(16#8A#, 8);
  gmul2_7(69) <= to_unsigned(16#8C#, 8);
  gmul2_7(70) <= to_unsigned(16#8E#, 8);
  gmul2_7(71) <= to_unsigned(16#90#, 8);
  gmul2_7(72) <= to_unsigned(16#92#, 8);
  gmul2_7(73) <= to_unsigned(16#94#, 8);
  gmul2_7(74) <= to_unsigned(16#96#, 8);
  gmul2_7(75) <= to_unsigned(16#98#, 8);
  gmul2_7(76) <= to_unsigned(16#9A#, 8);
  gmul2_7(77) <= to_unsigned(16#9C#, 8);
  gmul2_7(78) <= to_unsigned(16#9E#, 8);
  gmul2_7(79) <= to_unsigned(16#A0#, 8);
  gmul2_7(80) <= to_unsigned(16#A2#, 8);
  gmul2_7(81) <= to_unsigned(16#A4#, 8);
  gmul2_7(82) <= to_unsigned(16#A6#, 8);
  gmul2_7(83) <= to_unsigned(16#A8#, 8);
  gmul2_7(84) <= to_unsigned(16#AA#, 8);
  gmul2_7(85) <= to_unsigned(16#AC#, 8);
  gmul2_7(86) <= to_unsigned(16#AE#, 8);
  gmul2_7(87) <= to_unsigned(16#B0#, 8);
  gmul2_7(88) <= to_unsigned(16#B2#, 8);
  gmul2_7(89) <= to_unsigned(16#B4#, 8);
  gmul2_7(90) <= to_unsigned(16#B6#, 8);
  gmul2_7(91) <= to_unsigned(16#B8#, 8);
  gmul2_7(92) <= to_unsigned(16#BA#, 8);
  gmul2_7(93) <= to_unsigned(16#BC#, 8);
  gmul2_7(94) <= to_unsigned(16#BE#, 8);
  gmul2_7(95) <= to_unsigned(16#C0#, 8);
  gmul2_7(96) <= to_unsigned(16#C2#, 8);
  gmul2_7(97) <= to_unsigned(16#C4#, 8);
  gmul2_7(98) <= to_unsigned(16#C6#, 8);
  gmul2_7(99) <= to_unsigned(16#C8#, 8);
  gmul2_7(100) <= to_unsigned(16#CA#, 8);
  gmul2_7(101) <= to_unsigned(16#CC#, 8);
  gmul2_7(102) <= to_unsigned(16#CE#, 8);
  gmul2_7(103) <= to_unsigned(16#D0#, 8);
  gmul2_7(104) <= to_unsigned(16#D2#, 8);
  gmul2_7(105) <= to_unsigned(16#D4#, 8);
  gmul2_7(106) <= to_unsigned(16#D6#, 8);
  gmul2_7(107) <= to_unsigned(16#D8#, 8);
  gmul2_7(108) <= to_unsigned(16#DA#, 8);
  gmul2_7(109) <= to_unsigned(16#DC#, 8);
  gmul2_7(110) <= to_unsigned(16#DE#, 8);
  gmul2_7(111) <= to_unsigned(16#E0#, 8);
  gmul2_7(112) <= to_unsigned(16#E2#, 8);
  gmul2_7(113) <= to_unsigned(16#E4#, 8);
  gmul2_7(114) <= to_unsigned(16#E6#, 8);
  gmul2_7(115) <= to_unsigned(16#E8#, 8);
  gmul2_7(116) <= to_unsigned(16#EA#, 8);
  gmul2_7(117) <= to_unsigned(16#EC#, 8);
  gmul2_7(118) <= to_unsigned(16#EE#, 8);
  gmul2_7(119) <= to_unsigned(16#F0#, 8);
  gmul2_7(120) <= to_unsigned(16#F2#, 8);
  gmul2_7(121) <= to_unsigned(16#F4#, 8);
  gmul2_7(122) <= to_unsigned(16#F6#, 8);
  gmul2_7(123) <= to_unsigned(16#F8#, 8);
  gmul2_7(124) <= to_unsigned(16#FA#, 8);
  gmul2_7(125) <= to_unsigned(16#FC#, 8);
  gmul2_7(126) <= to_unsigned(16#FE#, 8);
  gmul2_7(127) <= to_unsigned(16#1B#, 8);
  gmul2_7(128) <= to_unsigned(16#19#, 8);
  gmul2_7(129) <= to_unsigned(16#1F#, 8);
  gmul2_7(130) <= to_unsigned(16#1D#, 8);
  gmul2_7(131) <= to_unsigned(16#13#, 8);
  gmul2_7(132) <= to_unsigned(16#11#, 8);
  gmul2_7(133) <= to_unsigned(16#17#, 8);
  gmul2_7(134) <= to_unsigned(16#15#, 8);
  gmul2_7(135) <= to_unsigned(16#0B#, 8);
  gmul2_7(136) <= to_unsigned(16#09#, 8);
  gmul2_7(137) <= to_unsigned(16#0F#, 8);
  gmul2_7(138) <= to_unsigned(16#0D#, 8);
  gmul2_7(139) <= to_unsigned(16#03#, 8);
  gmul2_7(140) <= to_unsigned(16#01#, 8);
  gmul2_7(141) <= to_unsigned(16#07#, 8);
  gmul2_7(142) <= to_unsigned(16#05#, 8);
  gmul2_7(143) <= to_unsigned(16#3B#, 8);
  gmul2_7(144) <= to_unsigned(16#39#, 8);
  gmul2_7(145) <= to_unsigned(16#3F#, 8);
  gmul2_7(146) <= to_unsigned(16#3D#, 8);
  gmul2_7(147) <= to_unsigned(16#33#, 8);
  gmul2_7(148) <= to_unsigned(16#31#, 8);
  gmul2_7(149) <= to_unsigned(16#37#, 8);
  gmul2_7(150) <= to_unsigned(16#35#, 8);
  gmul2_7(151) <= to_unsigned(16#2B#, 8);
  gmul2_7(152) <= to_unsigned(16#29#, 8);
  gmul2_7(153) <= to_unsigned(16#2F#, 8);
  gmul2_7(154) <= to_unsigned(16#2D#, 8);
  gmul2_7(155) <= to_unsigned(16#23#, 8);
  gmul2_7(156) <= to_unsigned(16#21#, 8);
  gmul2_7(157) <= to_unsigned(16#27#, 8);
  gmul2_7(158) <= to_unsigned(16#25#, 8);
  gmul2_7(159) <= to_unsigned(16#5B#, 8);
  gmul2_7(160) <= to_unsigned(16#59#, 8);
  gmul2_7(161) <= to_unsigned(16#5F#, 8);
  gmul2_7(162) <= to_unsigned(16#5D#, 8);
  gmul2_7(163) <= to_unsigned(16#53#, 8);
  gmul2_7(164) <= to_unsigned(16#51#, 8);
  gmul2_7(165) <= to_unsigned(16#57#, 8);
  gmul2_7(166) <= to_unsigned(16#55#, 8);
  gmul2_7(167) <= to_unsigned(16#4B#, 8);
  gmul2_7(168) <= to_unsigned(16#49#, 8);
  gmul2_7(169) <= to_unsigned(16#4F#, 8);
  gmul2_7(170) <= to_unsigned(16#4D#, 8);
  gmul2_7(171) <= to_unsigned(16#43#, 8);
  gmul2_7(172) <= to_unsigned(16#41#, 8);
  gmul2_7(173) <= to_unsigned(16#47#, 8);
  gmul2_7(174) <= to_unsigned(16#45#, 8);
  gmul2_7(175) <= to_unsigned(16#7B#, 8);
  gmul2_7(176) <= to_unsigned(16#79#, 8);
  gmul2_7(177) <= to_unsigned(16#7F#, 8);
  gmul2_7(178) <= to_unsigned(16#7D#, 8);
  gmul2_7(179) <= to_unsigned(16#73#, 8);
  gmul2_7(180) <= to_unsigned(16#71#, 8);
  gmul2_7(181) <= to_unsigned(16#77#, 8);
  gmul2_7(182) <= to_unsigned(16#75#, 8);
  gmul2_7(183) <= to_unsigned(16#6B#, 8);
  gmul2_7(184) <= to_unsigned(16#69#, 8);
  gmul2_7(185) <= to_unsigned(16#6F#, 8);
  gmul2_7(186) <= to_unsigned(16#6D#, 8);
  gmul2_7(187) <= to_unsigned(16#63#, 8);
  gmul2_7(188) <= to_unsigned(16#61#, 8);
  gmul2_7(189) <= to_unsigned(16#67#, 8);
  gmul2_7(190) <= to_unsigned(16#65#, 8);
  gmul2_7(191) <= to_unsigned(16#9B#, 8);
  gmul2_7(192) <= to_unsigned(16#99#, 8);
  gmul2_7(193) <= to_unsigned(16#9F#, 8);
  gmul2_7(194) <= to_unsigned(16#9D#, 8);
  gmul2_7(195) <= to_unsigned(16#93#, 8);
  gmul2_7(196) <= to_unsigned(16#91#, 8);
  gmul2_7(197) <= to_unsigned(16#97#, 8);
  gmul2_7(198) <= to_unsigned(16#95#, 8);
  gmul2_7(199) <= to_unsigned(16#8B#, 8);
  gmul2_7(200) <= to_unsigned(16#89#, 8);
  gmul2_7(201) <= to_unsigned(16#8F#, 8);
  gmul2_7(202) <= to_unsigned(16#8D#, 8);
  gmul2_7(203) <= to_unsigned(16#83#, 8);
  gmul2_7(204) <= to_unsigned(16#81#, 8);
  gmul2_7(205) <= to_unsigned(16#87#, 8);
  gmul2_7(206) <= to_unsigned(16#85#, 8);
  gmul2_7(207) <= to_unsigned(16#BB#, 8);
  gmul2_7(208) <= to_unsigned(16#B9#, 8);
  gmul2_7(209) <= to_unsigned(16#BF#, 8);
  gmul2_7(210) <= to_unsigned(16#BD#, 8);
  gmul2_7(211) <= to_unsigned(16#B3#, 8);
  gmul2_7(212) <= to_unsigned(16#B1#, 8);
  gmul2_7(213) <= to_unsigned(16#B7#, 8);
  gmul2_7(214) <= to_unsigned(16#B5#, 8);
  gmul2_7(215) <= to_unsigned(16#AB#, 8);
  gmul2_7(216) <= to_unsigned(16#A9#, 8);
  gmul2_7(217) <= to_unsigned(16#AF#, 8);
  gmul2_7(218) <= to_unsigned(16#AD#, 8);
  gmul2_7(219) <= to_unsigned(16#A3#, 8);
  gmul2_7(220) <= to_unsigned(16#A1#, 8);
  gmul2_7(221) <= to_unsigned(16#A7#, 8);
  gmul2_7(222) <= to_unsigned(16#A5#, 8);
  gmul2_7(223) <= to_unsigned(16#DB#, 8);
  gmul2_7(224) <= to_unsigned(16#D9#, 8);
  gmul2_7(225) <= to_unsigned(16#DF#, 8);
  gmul2_7(226) <= to_unsigned(16#DD#, 8);
  gmul2_7(227) <= to_unsigned(16#D3#, 8);
  gmul2_7(228) <= to_unsigned(16#D1#, 8);
  gmul2_7(229) <= to_unsigned(16#D7#, 8);
  gmul2_7(230) <= to_unsigned(16#D5#, 8);
  gmul2_7(231) <= to_unsigned(16#CB#, 8);
  gmul2_7(232) <= to_unsigned(16#C9#, 8);
  gmul2_7(233) <= to_unsigned(16#CF#, 8);
  gmul2_7(234) <= to_unsigned(16#CD#, 8);
  gmul2_7(235) <= to_unsigned(16#C3#, 8);
  gmul2_7(236) <= to_unsigned(16#C1#, 8);
  gmul2_7(237) <= to_unsigned(16#C7#, 8);
  gmul2_7(238) <= to_unsigned(16#C5#, 8);
  gmul2_7(239) <= to_unsigned(16#FB#, 8);
  gmul2_7(240) <= to_unsigned(16#F9#, 8);
  gmul2_7(241) <= to_unsigned(16#FF#, 8);
  gmul2_7(242) <= to_unsigned(16#FD#, 8);
  gmul2_7(243) <= to_unsigned(16#F3#, 8);
  gmul2_7(244) <= to_unsigned(16#F1#, 8);
  gmul2_7(245) <= to_unsigned(16#F7#, 8);
  gmul2_7(246) <= to_unsigned(16#F5#, 8);
  gmul2_7(247) <= to_unsigned(16#EB#, 8);
  gmul2_7(248) <= to_unsigned(16#E9#, 8);
  gmul2_7(249) <= to_unsigned(16#EF#, 8);
  gmul2_7(250) <= to_unsigned(16#ED#, 8);
  gmul2_7(251) <= to_unsigned(16#E3#, 8);
  gmul2_7(252) <= to_unsigned(16#E1#, 8);
  gmul2_7(253) <= to_unsigned(16#E7#, 8);
  gmul2_7(254) <= to_unsigned(16#E5#, 8);
  gmul2_7(255) <= to_unsigned(16#E5#, 8);

  gmul2_8(0) <= to_unsigned(16#02#, 8);
  gmul2_8(1) <= to_unsigned(16#04#, 8);
  gmul2_8(2) <= to_unsigned(16#06#, 8);
  gmul2_8(3) <= to_unsigned(16#08#, 8);
  gmul2_8(4) <= to_unsigned(16#0A#, 8);
  gmul2_8(5) <= to_unsigned(16#0C#, 8);
  gmul2_8(6) <= to_unsigned(16#0E#, 8);
  gmul2_8(7) <= to_unsigned(16#10#, 8);
  gmul2_8(8) <= to_unsigned(16#12#, 8);
  gmul2_8(9) <= to_unsigned(16#14#, 8);
  gmul2_8(10) <= to_unsigned(16#16#, 8);
  gmul2_8(11) <= to_unsigned(16#18#, 8);
  gmul2_8(12) <= to_unsigned(16#1A#, 8);
  gmul2_8(13) <= to_unsigned(16#1C#, 8);
  gmul2_8(14) <= to_unsigned(16#1E#, 8);
  gmul2_8(15) <= to_unsigned(16#20#, 8);
  gmul2_8(16) <= to_unsigned(16#22#, 8);
  gmul2_8(17) <= to_unsigned(16#24#, 8);
  gmul2_8(18) <= to_unsigned(16#26#, 8);
  gmul2_8(19) <= to_unsigned(16#28#, 8);
  gmul2_8(20) <= to_unsigned(16#2A#, 8);
  gmul2_8(21) <= to_unsigned(16#2C#, 8);
  gmul2_8(22) <= to_unsigned(16#2E#, 8);
  gmul2_8(23) <= to_unsigned(16#30#, 8);
  gmul2_8(24) <= to_unsigned(16#32#, 8);
  gmul2_8(25) <= to_unsigned(16#34#, 8);
  gmul2_8(26) <= to_unsigned(16#36#, 8);
  gmul2_8(27) <= to_unsigned(16#38#, 8);
  gmul2_8(28) <= to_unsigned(16#3A#, 8);
  gmul2_8(29) <= to_unsigned(16#3C#, 8);
  gmul2_8(30) <= to_unsigned(16#3E#, 8);
  gmul2_8(31) <= to_unsigned(16#40#, 8);
  gmul2_8(32) <= to_unsigned(16#42#, 8);
  gmul2_8(33) <= to_unsigned(16#44#, 8);
  gmul2_8(34) <= to_unsigned(16#46#, 8);
  gmul2_8(35) <= to_unsigned(16#48#, 8);
  gmul2_8(36) <= to_unsigned(16#4A#, 8);
  gmul2_8(37) <= to_unsigned(16#4C#, 8);
  gmul2_8(38) <= to_unsigned(16#4E#, 8);
  gmul2_8(39) <= to_unsigned(16#50#, 8);
  gmul2_8(40) <= to_unsigned(16#52#, 8);
  gmul2_8(41) <= to_unsigned(16#54#, 8);
  gmul2_8(42) <= to_unsigned(16#56#, 8);
  gmul2_8(43) <= to_unsigned(16#58#, 8);
  gmul2_8(44) <= to_unsigned(16#5A#, 8);
  gmul2_8(45) <= to_unsigned(16#5C#, 8);
  gmul2_8(46) <= to_unsigned(16#5E#, 8);
  gmul2_8(47) <= to_unsigned(16#60#, 8);
  gmul2_8(48) <= to_unsigned(16#62#, 8);
  gmul2_8(49) <= to_unsigned(16#64#, 8);
  gmul2_8(50) <= to_unsigned(16#66#, 8);
  gmul2_8(51) <= to_unsigned(16#68#, 8);
  gmul2_8(52) <= to_unsigned(16#6A#, 8);
  gmul2_8(53) <= to_unsigned(16#6C#, 8);
  gmul2_8(54) <= to_unsigned(16#6E#, 8);
  gmul2_8(55) <= to_unsigned(16#70#, 8);
  gmul2_8(56) <= to_unsigned(16#72#, 8);
  gmul2_8(57) <= to_unsigned(16#74#, 8);
  gmul2_8(58) <= to_unsigned(16#76#, 8);
  gmul2_8(59) <= to_unsigned(16#78#, 8);
  gmul2_8(60) <= to_unsigned(16#7A#, 8);
  gmul2_8(61) <= to_unsigned(16#7C#, 8);
  gmul2_8(62) <= to_unsigned(16#7E#, 8);
  gmul2_8(63) <= to_unsigned(16#80#, 8);
  gmul2_8(64) <= to_unsigned(16#82#, 8);
  gmul2_8(65) <= to_unsigned(16#84#, 8);
  gmul2_8(66) <= to_unsigned(16#86#, 8);
  gmul2_8(67) <= to_unsigned(16#88#, 8);
  gmul2_8(68) <= to_unsigned(16#8A#, 8);
  gmul2_8(69) <= to_unsigned(16#8C#, 8);
  gmul2_8(70) <= to_unsigned(16#8E#, 8);
  gmul2_8(71) <= to_unsigned(16#90#, 8);
  gmul2_8(72) <= to_unsigned(16#92#, 8);
  gmul2_8(73) <= to_unsigned(16#94#, 8);
  gmul2_8(74) <= to_unsigned(16#96#, 8);
  gmul2_8(75) <= to_unsigned(16#98#, 8);
  gmul2_8(76) <= to_unsigned(16#9A#, 8);
  gmul2_8(77) <= to_unsigned(16#9C#, 8);
  gmul2_8(78) <= to_unsigned(16#9E#, 8);
  gmul2_8(79) <= to_unsigned(16#A0#, 8);
  gmul2_8(80) <= to_unsigned(16#A2#, 8);
  gmul2_8(81) <= to_unsigned(16#A4#, 8);
  gmul2_8(82) <= to_unsigned(16#A6#, 8);
  gmul2_8(83) <= to_unsigned(16#A8#, 8);
  gmul2_8(84) <= to_unsigned(16#AA#, 8);
  gmul2_8(85) <= to_unsigned(16#AC#, 8);
  gmul2_8(86) <= to_unsigned(16#AE#, 8);
  gmul2_8(87) <= to_unsigned(16#B0#, 8);
  gmul2_8(88) <= to_unsigned(16#B2#, 8);
  gmul2_8(89) <= to_unsigned(16#B4#, 8);
  gmul2_8(90) <= to_unsigned(16#B6#, 8);
  gmul2_8(91) <= to_unsigned(16#B8#, 8);
  gmul2_8(92) <= to_unsigned(16#BA#, 8);
  gmul2_8(93) <= to_unsigned(16#BC#, 8);
  gmul2_8(94) <= to_unsigned(16#BE#, 8);
  gmul2_8(95) <= to_unsigned(16#C0#, 8);
  gmul2_8(96) <= to_unsigned(16#C2#, 8);
  gmul2_8(97) <= to_unsigned(16#C4#, 8);
  gmul2_8(98) <= to_unsigned(16#C6#, 8);
  gmul2_8(99) <= to_unsigned(16#C8#, 8);
  gmul2_8(100) <= to_unsigned(16#CA#, 8);
  gmul2_8(101) <= to_unsigned(16#CC#, 8);
  gmul2_8(102) <= to_unsigned(16#CE#, 8);
  gmul2_8(103) <= to_unsigned(16#D0#, 8);
  gmul2_8(104) <= to_unsigned(16#D2#, 8);
  gmul2_8(105) <= to_unsigned(16#D4#, 8);
  gmul2_8(106) <= to_unsigned(16#D6#, 8);
  gmul2_8(107) <= to_unsigned(16#D8#, 8);
  gmul2_8(108) <= to_unsigned(16#DA#, 8);
  gmul2_8(109) <= to_unsigned(16#DC#, 8);
  gmul2_8(110) <= to_unsigned(16#DE#, 8);
  gmul2_8(111) <= to_unsigned(16#E0#, 8);
  gmul2_8(112) <= to_unsigned(16#E2#, 8);
  gmul2_8(113) <= to_unsigned(16#E4#, 8);
  gmul2_8(114) <= to_unsigned(16#E6#, 8);
  gmul2_8(115) <= to_unsigned(16#E8#, 8);
  gmul2_8(116) <= to_unsigned(16#EA#, 8);
  gmul2_8(117) <= to_unsigned(16#EC#, 8);
  gmul2_8(118) <= to_unsigned(16#EE#, 8);
  gmul2_8(119) <= to_unsigned(16#F0#, 8);
  gmul2_8(120) <= to_unsigned(16#F2#, 8);
  gmul2_8(121) <= to_unsigned(16#F4#, 8);
  gmul2_8(122) <= to_unsigned(16#F6#, 8);
  gmul2_8(123) <= to_unsigned(16#F8#, 8);
  gmul2_8(124) <= to_unsigned(16#FA#, 8);
  gmul2_8(125) <= to_unsigned(16#FC#, 8);
  gmul2_8(126) <= to_unsigned(16#FE#, 8);
  gmul2_8(127) <= to_unsigned(16#1B#, 8);
  gmul2_8(128) <= to_unsigned(16#19#, 8);
  gmul2_8(129) <= to_unsigned(16#1F#, 8);
  gmul2_8(130) <= to_unsigned(16#1D#, 8);
  gmul2_8(131) <= to_unsigned(16#13#, 8);
  gmul2_8(132) <= to_unsigned(16#11#, 8);
  gmul2_8(133) <= to_unsigned(16#17#, 8);
  gmul2_8(134) <= to_unsigned(16#15#, 8);
  gmul2_8(135) <= to_unsigned(16#0B#, 8);
  gmul2_8(136) <= to_unsigned(16#09#, 8);
  gmul2_8(137) <= to_unsigned(16#0F#, 8);
  gmul2_8(138) <= to_unsigned(16#0D#, 8);
  gmul2_8(139) <= to_unsigned(16#03#, 8);
  gmul2_8(140) <= to_unsigned(16#01#, 8);
  gmul2_8(141) <= to_unsigned(16#07#, 8);
  gmul2_8(142) <= to_unsigned(16#05#, 8);
  gmul2_8(143) <= to_unsigned(16#3B#, 8);
  gmul2_8(144) <= to_unsigned(16#39#, 8);
  gmul2_8(145) <= to_unsigned(16#3F#, 8);
  gmul2_8(146) <= to_unsigned(16#3D#, 8);
  gmul2_8(147) <= to_unsigned(16#33#, 8);
  gmul2_8(148) <= to_unsigned(16#31#, 8);
  gmul2_8(149) <= to_unsigned(16#37#, 8);
  gmul2_8(150) <= to_unsigned(16#35#, 8);
  gmul2_8(151) <= to_unsigned(16#2B#, 8);
  gmul2_8(152) <= to_unsigned(16#29#, 8);
  gmul2_8(153) <= to_unsigned(16#2F#, 8);
  gmul2_8(154) <= to_unsigned(16#2D#, 8);
  gmul2_8(155) <= to_unsigned(16#23#, 8);
  gmul2_8(156) <= to_unsigned(16#21#, 8);
  gmul2_8(157) <= to_unsigned(16#27#, 8);
  gmul2_8(158) <= to_unsigned(16#25#, 8);
  gmul2_8(159) <= to_unsigned(16#5B#, 8);
  gmul2_8(160) <= to_unsigned(16#59#, 8);
  gmul2_8(161) <= to_unsigned(16#5F#, 8);
  gmul2_8(162) <= to_unsigned(16#5D#, 8);
  gmul2_8(163) <= to_unsigned(16#53#, 8);
  gmul2_8(164) <= to_unsigned(16#51#, 8);
  gmul2_8(165) <= to_unsigned(16#57#, 8);
  gmul2_8(166) <= to_unsigned(16#55#, 8);
  gmul2_8(167) <= to_unsigned(16#4B#, 8);
  gmul2_8(168) <= to_unsigned(16#49#, 8);
  gmul2_8(169) <= to_unsigned(16#4F#, 8);
  gmul2_8(170) <= to_unsigned(16#4D#, 8);
  gmul2_8(171) <= to_unsigned(16#43#, 8);
  gmul2_8(172) <= to_unsigned(16#41#, 8);
  gmul2_8(173) <= to_unsigned(16#47#, 8);
  gmul2_8(174) <= to_unsigned(16#45#, 8);
  gmul2_8(175) <= to_unsigned(16#7B#, 8);
  gmul2_8(176) <= to_unsigned(16#79#, 8);
  gmul2_8(177) <= to_unsigned(16#7F#, 8);
  gmul2_8(178) <= to_unsigned(16#7D#, 8);
  gmul2_8(179) <= to_unsigned(16#73#, 8);
  gmul2_8(180) <= to_unsigned(16#71#, 8);
  gmul2_8(181) <= to_unsigned(16#77#, 8);
  gmul2_8(182) <= to_unsigned(16#75#, 8);
  gmul2_8(183) <= to_unsigned(16#6B#, 8);
  gmul2_8(184) <= to_unsigned(16#69#, 8);
  gmul2_8(185) <= to_unsigned(16#6F#, 8);
  gmul2_8(186) <= to_unsigned(16#6D#, 8);
  gmul2_8(187) <= to_unsigned(16#63#, 8);
  gmul2_8(188) <= to_unsigned(16#61#, 8);
  gmul2_8(189) <= to_unsigned(16#67#, 8);
  gmul2_8(190) <= to_unsigned(16#65#, 8);
  gmul2_8(191) <= to_unsigned(16#9B#, 8);
  gmul2_8(192) <= to_unsigned(16#99#, 8);
  gmul2_8(193) <= to_unsigned(16#9F#, 8);
  gmul2_8(194) <= to_unsigned(16#9D#, 8);
  gmul2_8(195) <= to_unsigned(16#93#, 8);
  gmul2_8(196) <= to_unsigned(16#91#, 8);
  gmul2_8(197) <= to_unsigned(16#97#, 8);
  gmul2_8(198) <= to_unsigned(16#95#, 8);
  gmul2_8(199) <= to_unsigned(16#8B#, 8);
  gmul2_8(200) <= to_unsigned(16#89#, 8);
  gmul2_8(201) <= to_unsigned(16#8F#, 8);
  gmul2_8(202) <= to_unsigned(16#8D#, 8);
  gmul2_8(203) <= to_unsigned(16#83#, 8);
  gmul2_8(204) <= to_unsigned(16#81#, 8);
  gmul2_8(205) <= to_unsigned(16#87#, 8);
  gmul2_8(206) <= to_unsigned(16#85#, 8);
  gmul2_8(207) <= to_unsigned(16#BB#, 8);
  gmul2_8(208) <= to_unsigned(16#B9#, 8);
  gmul2_8(209) <= to_unsigned(16#BF#, 8);
  gmul2_8(210) <= to_unsigned(16#BD#, 8);
  gmul2_8(211) <= to_unsigned(16#B3#, 8);
  gmul2_8(212) <= to_unsigned(16#B1#, 8);
  gmul2_8(213) <= to_unsigned(16#B7#, 8);
  gmul2_8(214) <= to_unsigned(16#B5#, 8);
  gmul2_8(215) <= to_unsigned(16#AB#, 8);
  gmul2_8(216) <= to_unsigned(16#A9#, 8);
  gmul2_8(217) <= to_unsigned(16#AF#, 8);
  gmul2_8(218) <= to_unsigned(16#AD#, 8);
  gmul2_8(219) <= to_unsigned(16#A3#, 8);
  gmul2_8(220) <= to_unsigned(16#A1#, 8);
  gmul2_8(221) <= to_unsigned(16#A7#, 8);
  gmul2_8(222) <= to_unsigned(16#A5#, 8);
  gmul2_8(223) <= to_unsigned(16#DB#, 8);
  gmul2_8(224) <= to_unsigned(16#D9#, 8);
  gmul2_8(225) <= to_unsigned(16#DF#, 8);
  gmul2_8(226) <= to_unsigned(16#DD#, 8);
  gmul2_8(227) <= to_unsigned(16#D3#, 8);
  gmul2_8(228) <= to_unsigned(16#D1#, 8);
  gmul2_8(229) <= to_unsigned(16#D7#, 8);
  gmul2_8(230) <= to_unsigned(16#D5#, 8);
  gmul2_8(231) <= to_unsigned(16#CB#, 8);
  gmul2_8(232) <= to_unsigned(16#C9#, 8);
  gmul2_8(233) <= to_unsigned(16#CF#, 8);
  gmul2_8(234) <= to_unsigned(16#CD#, 8);
  gmul2_8(235) <= to_unsigned(16#C3#, 8);
  gmul2_8(236) <= to_unsigned(16#C1#, 8);
  gmul2_8(237) <= to_unsigned(16#C7#, 8);
  gmul2_8(238) <= to_unsigned(16#C5#, 8);
  gmul2_8(239) <= to_unsigned(16#FB#, 8);
  gmul2_8(240) <= to_unsigned(16#F9#, 8);
  gmul2_8(241) <= to_unsigned(16#FF#, 8);
  gmul2_8(242) <= to_unsigned(16#FD#, 8);
  gmul2_8(243) <= to_unsigned(16#F3#, 8);
  gmul2_8(244) <= to_unsigned(16#F1#, 8);
  gmul2_8(245) <= to_unsigned(16#F7#, 8);
  gmul2_8(246) <= to_unsigned(16#F5#, 8);
  gmul2_8(247) <= to_unsigned(16#EB#, 8);
  gmul2_8(248) <= to_unsigned(16#E9#, 8);
  gmul2_8(249) <= to_unsigned(16#EF#, 8);
  gmul2_8(250) <= to_unsigned(16#ED#, 8);
  gmul2_8(251) <= to_unsigned(16#E3#, 8);
  gmul2_8(252) <= to_unsigned(16#E1#, 8);
  gmul2_8(253) <= to_unsigned(16#E7#, 8);
  gmul2_8(254) <= to_unsigned(16#E5#, 8);
  gmul2_8(255) <= to_unsigned(16#E5#, 8);

  gmul3_8(0) <= to_unsigned(16#03#, 8);
  gmul3_8(1) <= to_unsigned(16#06#, 8);
  gmul3_8(2) <= to_unsigned(16#05#, 8);
  gmul3_8(3) <= to_unsigned(16#0C#, 8);
  gmul3_8(4) <= to_unsigned(16#0F#, 8);
  gmul3_8(5) <= to_unsigned(16#0A#, 8);
  gmul3_8(6) <= to_unsigned(16#09#, 8);
  gmul3_8(7) <= to_unsigned(16#18#, 8);
  gmul3_8(8) <= to_unsigned(16#1B#, 8);
  gmul3_8(9) <= to_unsigned(16#1E#, 8);
  gmul3_8(10) <= to_unsigned(16#1D#, 8);
  gmul3_8(11) <= to_unsigned(16#14#, 8);
  gmul3_8(12) <= to_unsigned(16#17#, 8);
  gmul3_8(13) <= to_unsigned(16#12#, 8);
  gmul3_8(14) <= to_unsigned(16#11#, 8);
  gmul3_8(15) <= to_unsigned(16#30#, 8);
  gmul3_8(16) <= to_unsigned(16#33#, 8);
  gmul3_8(17) <= to_unsigned(16#36#, 8);
  gmul3_8(18) <= to_unsigned(16#35#, 8);
  gmul3_8(19) <= to_unsigned(16#3C#, 8);
  gmul3_8(20) <= to_unsigned(16#3F#, 8);
  gmul3_8(21) <= to_unsigned(16#3A#, 8);
  gmul3_8(22) <= to_unsigned(16#39#, 8);
  gmul3_8(23) <= to_unsigned(16#28#, 8);
  gmul3_8(24) <= to_unsigned(16#2B#, 8);
  gmul3_8(25) <= to_unsigned(16#2E#, 8);
  gmul3_8(26) <= to_unsigned(16#2D#, 8);
  gmul3_8(27) <= to_unsigned(16#24#, 8);
  gmul3_8(28) <= to_unsigned(16#27#, 8);
  gmul3_8(29) <= to_unsigned(16#22#, 8);
  gmul3_8(30) <= to_unsigned(16#21#, 8);
  gmul3_8(31) <= to_unsigned(16#60#, 8);
  gmul3_8(32) <= to_unsigned(16#63#, 8);
  gmul3_8(33) <= to_unsigned(16#66#, 8);
  gmul3_8(34) <= to_unsigned(16#65#, 8);
  gmul3_8(35) <= to_unsigned(16#6C#, 8);
  gmul3_8(36) <= to_unsigned(16#6F#, 8);
  gmul3_8(37) <= to_unsigned(16#6A#, 8);
  gmul3_8(38) <= to_unsigned(16#69#, 8);
  gmul3_8(39) <= to_unsigned(16#78#, 8);
  gmul3_8(40) <= to_unsigned(16#7B#, 8);
  gmul3_8(41) <= to_unsigned(16#7E#, 8);
  gmul3_8(42) <= to_unsigned(16#7D#, 8);
  gmul3_8(43) <= to_unsigned(16#74#, 8);
  gmul3_8(44) <= to_unsigned(16#77#, 8);
  gmul3_8(45) <= to_unsigned(16#72#, 8);
  gmul3_8(46) <= to_unsigned(16#71#, 8);
  gmul3_8(47) <= to_unsigned(16#50#, 8);
  gmul3_8(48) <= to_unsigned(16#53#, 8);
  gmul3_8(49) <= to_unsigned(16#56#, 8);
  gmul3_8(50) <= to_unsigned(16#55#, 8);
  gmul3_8(51) <= to_unsigned(16#5C#, 8);
  gmul3_8(52) <= to_unsigned(16#5F#, 8);
  gmul3_8(53) <= to_unsigned(16#5A#, 8);
  gmul3_8(54) <= to_unsigned(16#59#, 8);
  gmul3_8(55) <= to_unsigned(16#48#, 8);
  gmul3_8(56) <= to_unsigned(16#4B#, 8);
  gmul3_8(57) <= to_unsigned(16#4E#, 8);
  gmul3_8(58) <= to_unsigned(16#4D#, 8);
  gmul3_8(59) <= to_unsigned(16#44#, 8);
  gmul3_8(60) <= to_unsigned(16#47#, 8);
  gmul3_8(61) <= to_unsigned(16#42#, 8);
  gmul3_8(62) <= to_unsigned(16#41#, 8);
  gmul3_8(63) <= to_unsigned(16#C0#, 8);
  gmul3_8(64) <= to_unsigned(16#C3#, 8);
  gmul3_8(65) <= to_unsigned(16#C6#, 8);
  gmul3_8(66) <= to_unsigned(16#C5#, 8);
  gmul3_8(67) <= to_unsigned(16#CC#, 8);
  gmul3_8(68) <= to_unsigned(16#CF#, 8);
  gmul3_8(69) <= to_unsigned(16#CA#, 8);
  gmul3_8(70) <= to_unsigned(16#C9#, 8);
  gmul3_8(71) <= to_unsigned(16#D8#, 8);
  gmul3_8(72) <= to_unsigned(16#DB#, 8);
  gmul3_8(73) <= to_unsigned(16#DE#, 8);
  gmul3_8(74) <= to_unsigned(16#DD#, 8);
  gmul3_8(75) <= to_unsigned(16#D4#, 8);
  gmul3_8(76) <= to_unsigned(16#D7#, 8);
  gmul3_8(77) <= to_unsigned(16#D2#, 8);
  gmul3_8(78) <= to_unsigned(16#D1#, 8);
  gmul3_8(79) <= to_unsigned(16#F0#, 8);
  gmul3_8(80) <= to_unsigned(16#F3#, 8);
  gmul3_8(81) <= to_unsigned(16#F6#, 8);
  gmul3_8(82) <= to_unsigned(16#F5#, 8);
  gmul3_8(83) <= to_unsigned(16#FC#, 8);
  gmul3_8(84) <= to_unsigned(16#FF#, 8);
  gmul3_8(85) <= to_unsigned(16#FA#, 8);
  gmul3_8(86) <= to_unsigned(16#F9#, 8);
  gmul3_8(87) <= to_unsigned(16#E8#, 8);
  gmul3_8(88) <= to_unsigned(16#EB#, 8);
  gmul3_8(89) <= to_unsigned(16#EE#, 8);
  gmul3_8(90) <= to_unsigned(16#ED#, 8);
  gmul3_8(91) <= to_unsigned(16#E4#, 8);
  gmul3_8(92) <= to_unsigned(16#E7#, 8);
  gmul3_8(93) <= to_unsigned(16#E2#, 8);
  gmul3_8(94) <= to_unsigned(16#E1#, 8);
  gmul3_8(95) <= to_unsigned(16#A0#, 8);
  gmul3_8(96) <= to_unsigned(16#A3#, 8);
  gmul3_8(97) <= to_unsigned(16#A6#, 8);
  gmul3_8(98) <= to_unsigned(16#A5#, 8);
  gmul3_8(99) <= to_unsigned(16#AC#, 8);
  gmul3_8(100) <= to_unsigned(16#AF#, 8);
  gmul3_8(101) <= to_unsigned(16#AA#, 8);
  gmul3_8(102) <= to_unsigned(16#A9#, 8);
  gmul3_8(103) <= to_unsigned(16#B8#, 8);
  gmul3_8(104) <= to_unsigned(16#BB#, 8);
  gmul3_8(105) <= to_unsigned(16#BE#, 8);
  gmul3_8(106) <= to_unsigned(16#BD#, 8);
  gmul3_8(107) <= to_unsigned(16#B4#, 8);
  gmul3_8(108) <= to_unsigned(16#B7#, 8);
  gmul3_8(109) <= to_unsigned(16#B2#, 8);
  gmul3_8(110) <= to_unsigned(16#B1#, 8);
  gmul3_8(111) <= to_unsigned(16#90#, 8);
  gmul3_8(112) <= to_unsigned(16#93#, 8);
  gmul3_8(113) <= to_unsigned(16#96#, 8);
  gmul3_8(114) <= to_unsigned(16#95#, 8);
  gmul3_8(115) <= to_unsigned(16#9C#, 8);
  gmul3_8(116) <= to_unsigned(16#9F#, 8);
  gmul3_8(117) <= to_unsigned(16#9A#, 8);
  gmul3_8(118) <= to_unsigned(16#99#, 8);
  gmul3_8(119) <= to_unsigned(16#88#, 8);
  gmul3_8(120) <= to_unsigned(16#8B#, 8);
  gmul3_8(121) <= to_unsigned(16#8E#, 8);
  gmul3_8(122) <= to_unsigned(16#8D#, 8);
  gmul3_8(123) <= to_unsigned(16#84#, 8);
  gmul3_8(124) <= to_unsigned(16#87#, 8);
  gmul3_8(125) <= to_unsigned(16#82#, 8);
  gmul3_8(126) <= to_unsigned(16#81#, 8);
  gmul3_8(127) <= to_unsigned(16#9B#, 8);
  gmul3_8(128) <= to_unsigned(16#98#, 8);
  gmul3_8(129) <= to_unsigned(16#9D#, 8);
  gmul3_8(130) <= to_unsigned(16#9E#, 8);
  gmul3_8(131) <= to_unsigned(16#97#, 8);
  gmul3_8(132) <= to_unsigned(16#94#, 8);
  gmul3_8(133) <= to_unsigned(16#91#, 8);
  gmul3_8(134) <= to_unsigned(16#92#, 8);
  gmul3_8(135) <= to_unsigned(16#83#, 8);
  gmul3_8(136) <= to_unsigned(16#80#, 8);
  gmul3_8(137) <= to_unsigned(16#85#, 8);
  gmul3_8(138) <= to_unsigned(16#86#, 8);
  gmul3_8(139) <= to_unsigned(16#8F#, 8);
  gmul3_8(140) <= to_unsigned(16#8C#, 8);
  gmul3_8(141) <= to_unsigned(16#89#, 8);
  gmul3_8(142) <= to_unsigned(16#8A#, 8);
  gmul3_8(143) <= to_unsigned(16#AB#, 8);
  gmul3_8(144) <= to_unsigned(16#A8#, 8);
  gmul3_8(145) <= to_unsigned(16#AD#, 8);
  gmul3_8(146) <= to_unsigned(16#AE#, 8);
  gmul3_8(147) <= to_unsigned(16#A7#, 8);
  gmul3_8(148) <= to_unsigned(16#A4#, 8);
  gmul3_8(149) <= to_unsigned(16#A1#, 8);
  gmul3_8(150) <= to_unsigned(16#A2#, 8);
  gmul3_8(151) <= to_unsigned(16#B3#, 8);
  gmul3_8(152) <= to_unsigned(16#B0#, 8);
  gmul3_8(153) <= to_unsigned(16#B5#, 8);
  gmul3_8(154) <= to_unsigned(16#B6#, 8);
  gmul3_8(155) <= to_unsigned(16#BF#, 8);
  gmul3_8(156) <= to_unsigned(16#BC#, 8);
  gmul3_8(157) <= to_unsigned(16#B9#, 8);
  gmul3_8(158) <= to_unsigned(16#BA#, 8);
  gmul3_8(159) <= to_unsigned(16#FB#, 8);
  gmul3_8(160) <= to_unsigned(16#F8#, 8);
  gmul3_8(161) <= to_unsigned(16#FD#, 8);
  gmul3_8(162) <= to_unsigned(16#FE#, 8);
  gmul3_8(163) <= to_unsigned(16#F7#, 8);
  gmul3_8(164) <= to_unsigned(16#F4#, 8);
  gmul3_8(165) <= to_unsigned(16#F1#, 8);
  gmul3_8(166) <= to_unsigned(16#F2#, 8);
  gmul3_8(167) <= to_unsigned(16#E3#, 8);
  gmul3_8(168) <= to_unsigned(16#E0#, 8);
  gmul3_8(169) <= to_unsigned(16#E5#, 8);
  gmul3_8(170) <= to_unsigned(16#E6#, 8);
  gmul3_8(171) <= to_unsigned(16#EF#, 8);
  gmul3_8(172) <= to_unsigned(16#EC#, 8);
  gmul3_8(173) <= to_unsigned(16#E9#, 8);
  gmul3_8(174) <= to_unsigned(16#EA#, 8);
  gmul3_8(175) <= to_unsigned(16#CB#, 8);
  gmul3_8(176) <= to_unsigned(16#C8#, 8);
  gmul3_8(177) <= to_unsigned(16#CD#, 8);
  gmul3_8(178) <= to_unsigned(16#CE#, 8);
  gmul3_8(179) <= to_unsigned(16#C7#, 8);
  gmul3_8(180) <= to_unsigned(16#C4#, 8);
  gmul3_8(181) <= to_unsigned(16#C1#, 8);
  gmul3_8(182) <= to_unsigned(16#C2#, 8);
  gmul3_8(183) <= to_unsigned(16#D3#, 8);
  gmul3_8(184) <= to_unsigned(16#D0#, 8);
  gmul3_8(185) <= to_unsigned(16#D5#, 8);
  gmul3_8(186) <= to_unsigned(16#D6#, 8);
  gmul3_8(187) <= to_unsigned(16#DF#, 8);
  gmul3_8(188) <= to_unsigned(16#DC#, 8);
  gmul3_8(189) <= to_unsigned(16#D9#, 8);
  gmul3_8(190) <= to_unsigned(16#DA#, 8);
  gmul3_8(191) <= to_unsigned(16#5B#, 8);
  gmul3_8(192) <= to_unsigned(16#58#, 8);
  gmul3_8(193) <= to_unsigned(16#5D#, 8);
  gmul3_8(194) <= to_unsigned(16#5E#, 8);
  gmul3_8(195) <= to_unsigned(16#57#, 8);
  gmul3_8(196) <= to_unsigned(16#54#, 8);
  gmul3_8(197) <= to_unsigned(16#51#, 8);
  gmul3_8(198) <= to_unsigned(16#52#, 8);
  gmul3_8(199) <= to_unsigned(16#43#, 8);
  gmul3_8(200) <= to_unsigned(16#40#, 8);
  gmul3_8(201) <= to_unsigned(16#45#, 8);
  gmul3_8(202) <= to_unsigned(16#46#, 8);
  gmul3_8(203) <= to_unsigned(16#4F#, 8);
  gmul3_8(204) <= to_unsigned(16#4C#, 8);
  gmul3_8(205) <= to_unsigned(16#49#, 8);
  gmul3_8(206) <= to_unsigned(16#4A#, 8);
  gmul3_8(207) <= to_unsigned(16#6B#, 8);
  gmul3_8(208) <= to_unsigned(16#68#, 8);
  gmul3_8(209) <= to_unsigned(16#6D#, 8);
  gmul3_8(210) <= to_unsigned(16#6E#, 8);
  gmul3_8(211) <= to_unsigned(16#67#, 8);
  gmul3_8(212) <= to_unsigned(16#64#, 8);
  gmul3_8(213) <= to_unsigned(16#61#, 8);
  gmul3_8(214) <= to_unsigned(16#62#, 8);
  gmul3_8(215) <= to_unsigned(16#73#, 8);
  gmul3_8(216) <= to_unsigned(16#70#, 8);
  gmul3_8(217) <= to_unsigned(16#75#, 8);
  gmul3_8(218) <= to_unsigned(16#76#, 8);
  gmul3_8(219) <= to_unsigned(16#7F#, 8);
  gmul3_8(220) <= to_unsigned(16#7C#, 8);
  gmul3_8(221) <= to_unsigned(16#79#, 8);
  gmul3_8(222) <= to_unsigned(16#7A#, 8);
  gmul3_8(223) <= to_unsigned(16#3B#, 8);
  gmul3_8(224) <= to_unsigned(16#38#, 8);
  gmul3_8(225) <= to_unsigned(16#3D#, 8);
  gmul3_8(226) <= to_unsigned(16#3E#, 8);
  gmul3_8(227) <= to_unsigned(16#37#, 8);
  gmul3_8(228) <= to_unsigned(16#34#, 8);
  gmul3_8(229) <= to_unsigned(16#31#, 8);
  gmul3_8(230) <= to_unsigned(16#32#, 8);
  gmul3_8(231) <= to_unsigned(16#23#, 8);
  gmul3_8(232) <= to_unsigned(16#20#, 8);
  gmul3_8(233) <= to_unsigned(16#25#, 8);
  gmul3_8(234) <= to_unsigned(16#26#, 8);
  gmul3_8(235) <= to_unsigned(16#2F#, 8);
  gmul3_8(236) <= to_unsigned(16#2C#, 8);
  gmul3_8(237) <= to_unsigned(16#29#, 8);
  gmul3_8(238) <= to_unsigned(16#2A#, 8);
  gmul3_8(239) <= to_unsigned(16#0B#, 8);
  gmul3_8(240) <= to_unsigned(16#08#, 8);
  gmul3_8(241) <= to_unsigned(16#0D#, 8);
  gmul3_8(242) <= to_unsigned(16#0E#, 8);
  gmul3_8(243) <= to_unsigned(16#07#, 8);
  gmul3_8(244) <= to_unsigned(16#04#, 8);
  gmul3_8(245) <= to_unsigned(16#01#, 8);
  gmul3_8(246) <= to_unsigned(16#02#, 8);
  gmul3_8(247) <= to_unsigned(16#13#, 8);
  gmul3_8(248) <= to_unsigned(16#10#, 8);
  gmul3_8(249) <= to_unsigned(16#15#, 8);
  gmul3_8(250) <= to_unsigned(16#16#, 8);
  gmul3_8(251) <= to_unsigned(16#1F#, 8);
  gmul3_8(252) <= to_unsigned(16#1C#, 8);
  gmul3_8(253) <= to_unsigned(16#19#, 8);
  gmul3_8(254) <= to_unsigned(16#1A#, 8);
  gmul3_8(255) <= to_unsigned(16#1A#, 8);

  gmul2_9(0) <= to_unsigned(16#02#, 8);
  gmul2_9(1) <= to_unsigned(16#04#, 8);
  gmul2_9(2) <= to_unsigned(16#06#, 8);
  gmul2_9(3) <= to_unsigned(16#08#, 8);
  gmul2_9(4) <= to_unsigned(16#0A#, 8);
  gmul2_9(5) <= to_unsigned(16#0C#, 8);
  gmul2_9(6) <= to_unsigned(16#0E#, 8);
  gmul2_9(7) <= to_unsigned(16#10#, 8);
  gmul2_9(8) <= to_unsigned(16#12#, 8);
  gmul2_9(9) <= to_unsigned(16#14#, 8);
  gmul2_9(10) <= to_unsigned(16#16#, 8);
  gmul2_9(11) <= to_unsigned(16#18#, 8);
  gmul2_9(12) <= to_unsigned(16#1A#, 8);
  gmul2_9(13) <= to_unsigned(16#1C#, 8);
  gmul2_9(14) <= to_unsigned(16#1E#, 8);
  gmul2_9(15) <= to_unsigned(16#20#, 8);
  gmul2_9(16) <= to_unsigned(16#22#, 8);
  gmul2_9(17) <= to_unsigned(16#24#, 8);
  gmul2_9(18) <= to_unsigned(16#26#, 8);
  gmul2_9(19) <= to_unsigned(16#28#, 8);
  gmul2_9(20) <= to_unsigned(16#2A#, 8);
  gmul2_9(21) <= to_unsigned(16#2C#, 8);
  gmul2_9(22) <= to_unsigned(16#2E#, 8);
  gmul2_9(23) <= to_unsigned(16#30#, 8);
  gmul2_9(24) <= to_unsigned(16#32#, 8);
  gmul2_9(25) <= to_unsigned(16#34#, 8);
  gmul2_9(26) <= to_unsigned(16#36#, 8);
  gmul2_9(27) <= to_unsigned(16#38#, 8);
  gmul2_9(28) <= to_unsigned(16#3A#, 8);
  gmul2_9(29) <= to_unsigned(16#3C#, 8);
  gmul2_9(30) <= to_unsigned(16#3E#, 8);
  gmul2_9(31) <= to_unsigned(16#40#, 8);
  gmul2_9(32) <= to_unsigned(16#42#, 8);
  gmul2_9(33) <= to_unsigned(16#44#, 8);
  gmul2_9(34) <= to_unsigned(16#46#, 8);
  gmul2_9(35) <= to_unsigned(16#48#, 8);
  gmul2_9(36) <= to_unsigned(16#4A#, 8);
  gmul2_9(37) <= to_unsigned(16#4C#, 8);
  gmul2_9(38) <= to_unsigned(16#4E#, 8);
  gmul2_9(39) <= to_unsigned(16#50#, 8);
  gmul2_9(40) <= to_unsigned(16#52#, 8);
  gmul2_9(41) <= to_unsigned(16#54#, 8);
  gmul2_9(42) <= to_unsigned(16#56#, 8);
  gmul2_9(43) <= to_unsigned(16#58#, 8);
  gmul2_9(44) <= to_unsigned(16#5A#, 8);
  gmul2_9(45) <= to_unsigned(16#5C#, 8);
  gmul2_9(46) <= to_unsigned(16#5E#, 8);
  gmul2_9(47) <= to_unsigned(16#60#, 8);
  gmul2_9(48) <= to_unsigned(16#62#, 8);
  gmul2_9(49) <= to_unsigned(16#64#, 8);
  gmul2_9(50) <= to_unsigned(16#66#, 8);
  gmul2_9(51) <= to_unsigned(16#68#, 8);
  gmul2_9(52) <= to_unsigned(16#6A#, 8);
  gmul2_9(53) <= to_unsigned(16#6C#, 8);
  gmul2_9(54) <= to_unsigned(16#6E#, 8);
  gmul2_9(55) <= to_unsigned(16#70#, 8);
  gmul2_9(56) <= to_unsigned(16#72#, 8);
  gmul2_9(57) <= to_unsigned(16#74#, 8);
  gmul2_9(58) <= to_unsigned(16#76#, 8);
  gmul2_9(59) <= to_unsigned(16#78#, 8);
  gmul2_9(60) <= to_unsigned(16#7A#, 8);
  gmul2_9(61) <= to_unsigned(16#7C#, 8);
  gmul2_9(62) <= to_unsigned(16#7E#, 8);
  gmul2_9(63) <= to_unsigned(16#80#, 8);
  gmul2_9(64) <= to_unsigned(16#82#, 8);
  gmul2_9(65) <= to_unsigned(16#84#, 8);
  gmul2_9(66) <= to_unsigned(16#86#, 8);
  gmul2_9(67) <= to_unsigned(16#88#, 8);
  gmul2_9(68) <= to_unsigned(16#8A#, 8);
  gmul2_9(69) <= to_unsigned(16#8C#, 8);
  gmul2_9(70) <= to_unsigned(16#8E#, 8);
  gmul2_9(71) <= to_unsigned(16#90#, 8);
  gmul2_9(72) <= to_unsigned(16#92#, 8);
  gmul2_9(73) <= to_unsigned(16#94#, 8);
  gmul2_9(74) <= to_unsigned(16#96#, 8);
  gmul2_9(75) <= to_unsigned(16#98#, 8);
  gmul2_9(76) <= to_unsigned(16#9A#, 8);
  gmul2_9(77) <= to_unsigned(16#9C#, 8);
  gmul2_9(78) <= to_unsigned(16#9E#, 8);
  gmul2_9(79) <= to_unsigned(16#A0#, 8);
  gmul2_9(80) <= to_unsigned(16#A2#, 8);
  gmul2_9(81) <= to_unsigned(16#A4#, 8);
  gmul2_9(82) <= to_unsigned(16#A6#, 8);
  gmul2_9(83) <= to_unsigned(16#A8#, 8);
  gmul2_9(84) <= to_unsigned(16#AA#, 8);
  gmul2_9(85) <= to_unsigned(16#AC#, 8);
  gmul2_9(86) <= to_unsigned(16#AE#, 8);
  gmul2_9(87) <= to_unsigned(16#B0#, 8);
  gmul2_9(88) <= to_unsigned(16#B2#, 8);
  gmul2_9(89) <= to_unsigned(16#B4#, 8);
  gmul2_9(90) <= to_unsigned(16#B6#, 8);
  gmul2_9(91) <= to_unsigned(16#B8#, 8);
  gmul2_9(92) <= to_unsigned(16#BA#, 8);
  gmul2_9(93) <= to_unsigned(16#BC#, 8);
  gmul2_9(94) <= to_unsigned(16#BE#, 8);
  gmul2_9(95) <= to_unsigned(16#C0#, 8);
  gmul2_9(96) <= to_unsigned(16#C2#, 8);
  gmul2_9(97) <= to_unsigned(16#C4#, 8);
  gmul2_9(98) <= to_unsigned(16#C6#, 8);
  gmul2_9(99) <= to_unsigned(16#C8#, 8);
  gmul2_9(100) <= to_unsigned(16#CA#, 8);
  gmul2_9(101) <= to_unsigned(16#CC#, 8);
  gmul2_9(102) <= to_unsigned(16#CE#, 8);
  gmul2_9(103) <= to_unsigned(16#D0#, 8);
  gmul2_9(104) <= to_unsigned(16#D2#, 8);
  gmul2_9(105) <= to_unsigned(16#D4#, 8);
  gmul2_9(106) <= to_unsigned(16#D6#, 8);
  gmul2_9(107) <= to_unsigned(16#D8#, 8);
  gmul2_9(108) <= to_unsigned(16#DA#, 8);
  gmul2_9(109) <= to_unsigned(16#DC#, 8);
  gmul2_9(110) <= to_unsigned(16#DE#, 8);
  gmul2_9(111) <= to_unsigned(16#E0#, 8);
  gmul2_9(112) <= to_unsigned(16#E2#, 8);
  gmul2_9(113) <= to_unsigned(16#E4#, 8);
  gmul2_9(114) <= to_unsigned(16#E6#, 8);
  gmul2_9(115) <= to_unsigned(16#E8#, 8);
  gmul2_9(116) <= to_unsigned(16#EA#, 8);
  gmul2_9(117) <= to_unsigned(16#EC#, 8);
  gmul2_9(118) <= to_unsigned(16#EE#, 8);
  gmul2_9(119) <= to_unsigned(16#F0#, 8);
  gmul2_9(120) <= to_unsigned(16#F2#, 8);
  gmul2_9(121) <= to_unsigned(16#F4#, 8);
  gmul2_9(122) <= to_unsigned(16#F6#, 8);
  gmul2_9(123) <= to_unsigned(16#F8#, 8);
  gmul2_9(124) <= to_unsigned(16#FA#, 8);
  gmul2_9(125) <= to_unsigned(16#FC#, 8);
  gmul2_9(126) <= to_unsigned(16#FE#, 8);
  gmul2_9(127) <= to_unsigned(16#1B#, 8);
  gmul2_9(128) <= to_unsigned(16#19#, 8);
  gmul2_9(129) <= to_unsigned(16#1F#, 8);
  gmul2_9(130) <= to_unsigned(16#1D#, 8);
  gmul2_9(131) <= to_unsigned(16#13#, 8);
  gmul2_9(132) <= to_unsigned(16#11#, 8);
  gmul2_9(133) <= to_unsigned(16#17#, 8);
  gmul2_9(134) <= to_unsigned(16#15#, 8);
  gmul2_9(135) <= to_unsigned(16#0B#, 8);
  gmul2_9(136) <= to_unsigned(16#09#, 8);
  gmul2_9(137) <= to_unsigned(16#0F#, 8);
  gmul2_9(138) <= to_unsigned(16#0D#, 8);
  gmul2_9(139) <= to_unsigned(16#03#, 8);
  gmul2_9(140) <= to_unsigned(16#01#, 8);
  gmul2_9(141) <= to_unsigned(16#07#, 8);
  gmul2_9(142) <= to_unsigned(16#05#, 8);
  gmul2_9(143) <= to_unsigned(16#3B#, 8);
  gmul2_9(144) <= to_unsigned(16#39#, 8);
  gmul2_9(145) <= to_unsigned(16#3F#, 8);
  gmul2_9(146) <= to_unsigned(16#3D#, 8);
  gmul2_9(147) <= to_unsigned(16#33#, 8);
  gmul2_9(148) <= to_unsigned(16#31#, 8);
  gmul2_9(149) <= to_unsigned(16#37#, 8);
  gmul2_9(150) <= to_unsigned(16#35#, 8);
  gmul2_9(151) <= to_unsigned(16#2B#, 8);
  gmul2_9(152) <= to_unsigned(16#29#, 8);
  gmul2_9(153) <= to_unsigned(16#2F#, 8);
  gmul2_9(154) <= to_unsigned(16#2D#, 8);
  gmul2_9(155) <= to_unsigned(16#23#, 8);
  gmul2_9(156) <= to_unsigned(16#21#, 8);
  gmul2_9(157) <= to_unsigned(16#27#, 8);
  gmul2_9(158) <= to_unsigned(16#25#, 8);
  gmul2_9(159) <= to_unsigned(16#5B#, 8);
  gmul2_9(160) <= to_unsigned(16#59#, 8);
  gmul2_9(161) <= to_unsigned(16#5F#, 8);
  gmul2_9(162) <= to_unsigned(16#5D#, 8);
  gmul2_9(163) <= to_unsigned(16#53#, 8);
  gmul2_9(164) <= to_unsigned(16#51#, 8);
  gmul2_9(165) <= to_unsigned(16#57#, 8);
  gmul2_9(166) <= to_unsigned(16#55#, 8);
  gmul2_9(167) <= to_unsigned(16#4B#, 8);
  gmul2_9(168) <= to_unsigned(16#49#, 8);
  gmul2_9(169) <= to_unsigned(16#4F#, 8);
  gmul2_9(170) <= to_unsigned(16#4D#, 8);
  gmul2_9(171) <= to_unsigned(16#43#, 8);
  gmul2_9(172) <= to_unsigned(16#41#, 8);
  gmul2_9(173) <= to_unsigned(16#47#, 8);
  gmul2_9(174) <= to_unsigned(16#45#, 8);
  gmul2_9(175) <= to_unsigned(16#7B#, 8);
  gmul2_9(176) <= to_unsigned(16#79#, 8);
  gmul2_9(177) <= to_unsigned(16#7F#, 8);
  gmul2_9(178) <= to_unsigned(16#7D#, 8);
  gmul2_9(179) <= to_unsigned(16#73#, 8);
  gmul2_9(180) <= to_unsigned(16#71#, 8);
  gmul2_9(181) <= to_unsigned(16#77#, 8);
  gmul2_9(182) <= to_unsigned(16#75#, 8);
  gmul2_9(183) <= to_unsigned(16#6B#, 8);
  gmul2_9(184) <= to_unsigned(16#69#, 8);
  gmul2_9(185) <= to_unsigned(16#6F#, 8);
  gmul2_9(186) <= to_unsigned(16#6D#, 8);
  gmul2_9(187) <= to_unsigned(16#63#, 8);
  gmul2_9(188) <= to_unsigned(16#61#, 8);
  gmul2_9(189) <= to_unsigned(16#67#, 8);
  gmul2_9(190) <= to_unsigned(16#65#, 8);
  gmul2_9(191) <= to_unsigned(16#9B#, 8);
  gmul2_9(192) <= to_unsigned(16#99#, 8);
  gmul2_9(193) <= to_unsigned(16#9F#, 8);
  gmul2_9(194) <= to_unsigned(16#9D#, 8);
  gmul2_9(195) <= to_unsigned(16#93#, 8);
  gmul2_9(196) <= to_unsigned(16#91#, 8);
  gmul2_9(197) <= to_unsigned(16#97#, 8);
  gmul2_9(198) <= to_unsigned(16#95#, 8);
  gmul2_9(199) <= to_unsigned(16#8B#, 8);
  gmul2_9(200) <= to_unsigned(16#89#, 8);
  gmul2_9(201) <= to_unsigned(16#8F#, 8);
  gmul2_9(202) <= to_unsigned(16#8D#, 8);
  gmul2_9(203) <= to_unsigned(16#83#, 8);
  gmul2_9(204) <= to_unsigned(16#81#, 8);
  gmul2_9(205) <= to_unsigned(16#87#, 8);
  gmul2_9(206) <= to_unsigned(16#85#, 8);
  gmul2_9(207) <= to_unsigned(16#BB#, 8);
  gmul2_9(208) <= to_unsigned(16#B9#, 8);
  gmul2_9(209) <= to_unsigned(16#BF#, 8);
  gmul2_9(210) <= to_unsigned(16#BD#, 8);
  gmul2_9(211) <= to_unsigned(16#B3#, 8);
  gmul2_9(212) <= to_unsigned(16#B1#, 8);
  gmul2_9(213) <= to_unsigned(16#B7#, 8);
  gmul2_9(214) <= to_unsigned(16#B5#, 8);
  gmul2_9(215) <= to_unsigned(16#AB#, 8);
  gmul2_9(216) <= to_unsigned(16#A9#, 8);
  gmul2_9(217) <= to_unsigned(16#AF#, 8);
  gmul2_9(218) <= to_unsigned(16#AD#, 8);
  gmul2_9(219) <= to_unsigned(16#A3#, 8);
  gmul2_9(220) <= to_unsigned(16#A1#, 8);
  gmul2_9(221) <= to_unsigned(16#A7#, 8);
  gmul2_9(222) <= to_unsigned(16#A5#, 8);
  gmul2_9(223) <= to_unsigned(16#DB#, 8);
  gmul2_9(224) <= to_unsigned(16#D9#, 8);
  gmul2_9(225) <= to_unsigned(16#DF#, 8);
  gmul2_9(226) <= to_unsigned(16#DD#, 8);
  gmul2_9(227) <= to_unsigned(16#D3#, 8);
  gmul2_9(228) <= to_unsigned(16#D1#, 8);
  gmul2_9(229) <= to_unsigned(16#D7#, 8);
  gmul2_9(230) <= to_unsigned(16#D5#, 8);
  gmul2_9(231) <= to_unsigned(16#CB#, 8);
  gmul2_9(232) <= to_unsigned(16#C9#, 8);
  gmul2_9(233) <= to_unsigned(16#CF#, 8);
  gmul2_9(234) <= to_unsigned(16#CD#, 8);
  gmul2_9(235) <= to_unsigned(16#C3#, 8);
  gmul2_9(236) <= to_unsigned(16#C1#, 8);
  gmul2_9(237) <= to_unsigned(16#C7#, 8);
  gmul2_9(238) <= to_unsigned(16#C5#, 8);
  gmul2_9(239) <= to_unsigned(16#FB#, 8);
  gmul2_9(240) <= to_unsigned(16#F9#, 8);
  gmul2_9(241) <= to_unsigned(16#FF#, 8);
  gmul2_9(242) <= to_unsigned(16#FD#, 8);
  gmul2_9(243) <= to_unsigned(16#F3#, 8);
  gmul2_9(244) <= to_unsigned(16#F1#, 8);
  gmul2_9(245) <= to_unsigned(16#F7#, 8);
  gmul2_9(246) <= to_unsigned(16#F5#, 8);
  gmul2_9(247) <= to_unsigned(16#EB#, 8);
  gmul2_9(248) <= to_unsigned(16#E9#, 8);
  gmul2_9(249) <= to_unsigned(16#EF#, 8);
  gmul2_9(250) <= to_unsigned(16#ED#, 8);
  gmul2_9(251) <= to_unsigned(16#E3#, 8);
  gmul2_9(252) <= to_unsigned(16#E1#, 8);
  gmul2_9(253) <= to_unsigned(16#E7#, 8);
  gmul2_9(254) <= to_unsigned(16#E5#, 8);
  gmul2_9(255) <= to_unsigned(16#E5#, 8);

  gmul3_9(0) <= to_unsigned(16#03#, 8);
  gmul3_9(1) <= to_unsigned(16#06#, 8);
  gmul3_9(2) <= to_unsigned(16#05#, 8);
  gmul3_9(3) <= to_unsigned(16#0C#, 8);
  gmul3_9(4) <= to_unsigned(16#0F#, 8);
  gmul3_9(5) <= to_unsigned(16#0A#, 8);
  gmul3_9(6) <= to_unsigned(16#09#, 8);
  gmul3_9(7) <= to_unsigned(16#18#, 8);
  gmul3_9(8) <= to_unsigned(16#1B#, 8);
  gmul3_9(9) <= to_unsigned(16#1E#, 8);
  gmul3_9(10) <= to_unsigned(16#1D#, 8);
  gmul3_9(11) <= to_unsigned(16#14#, 8);
  gmul3_9(12) <= to_unsigned(16#17#, 8);
  gmul3_9(13) <= to_unsigned(16#12#, 8);
  gmul3_9(14) <= to_unsigned(16#11#, 8);
  gmul3_9(15) <= to_unsigned(16#30#, 8);
  gmul3_9(16) <= to_unsigned(16#33#, 8);
  gmul3_9(17) <= to_unsigned(16#36#, 8);
  gmul3_9(18) <= to_unsigned(16#35#, 8);
  gmul3_9(19) <= to_unsigned(16#3C#, 8);
  gmul3_9(20) <= to_unsigned(16#3F#, 8);
  gmul3_9(21) <= to_unsigned(16#3A#, 8);
  gmul3_9(22) <= to_unsigned(16#39#, 8);
  gmul3_9(23) <= to_unsigned(16#28#, 8);
  gmul3_9(24) <= to_unsigned(16#2B#, 8);
  gmul3_9(25) <= to_unsigned(16#2E#, 8);
  gmul3_9(26) <= to_unsigned(16#2D#, 8);
  gmul3_9(27) <= to_unsigned(16#24#, 8);
  gmul3_9(28) <= to_unsigned(16#27#, 8);
  gmul3_9(29) <= to_unsigned(16#22#, 8);
  gmul3_9(30) <= to_unsigned(16#21#, 8);
  gmul3_9(31) <= to_unsigned(16#60#, 8);
  gmul3_9(32) <= to_unsigned(16#63#, 8);
  gmul3_9(33) <= to_unsigned(16#66#, 8);
  gmul3_9(34) <= to_unsigned(16#65#, 8);
  gmul3_9(35) <= to_unsigned(16#6C#, 8);
  gmul3_9(36) <= to_unsigned(16#6F#, 8);
  gmul3_9(37) <= to_unsigned(16#6A#, 8);
  gmul3_9(38) <= to_unsigned(16#69#, 8);
  gmul3_9(39) <= to_unsigned(16#78#, 8);
  gmul3_9(40) <= to_unsigned(16#7B#, 8);
  gmul3_9(41) <= to_unsigned(16#7E#, 8);
  gmul3_9(42) <= to_unsigned(16#7D#, 8);
  gmul3_9(43) <= to_unsigned(16#74#, 8);
  gmul3_9(44) <= to_unsigned(16#77#, 8);
  gmul3_9(45) <= to_unsigned(16#72#, 8);
  gmul3_9(46) <= to_unsigned(16#71#, 8);
  gmul3_9(47) <= to_unsigned(16#50#, 8);
  gmul3_9(48) <= to_unsigned(16#53#, 8);
  gmul3_9(49) <= to_unsigned(16#56#, 8);
  gmul3_9(50) <= to_unsigned(16#55#, 8);
  gmul3_9(51) <= to_unsigned(16#5C#, 8);
  gmul3_9(52) <= to_unsigned(16#5F#, 8);
  gmul3_9(53) <= to_unsigned(16#5A#, 8);
  gmul3_9(54) <= to_unsigned(16#59#, 8);
  gmul3_9(55) <= to_unsigned(16#48#, 8);
  gmul3_9(56) <= to_unsigned(16#4B#, 8);
  gmul3_9(57) <= to_unsigned(16#4E#, 8);
  gmul3_9(58) <= to_unsigned(16#4D#, 8);
  gmul3_9(59) <= to_unsigned(16#44#, 8);
  gmul3_9(60) <= to_unsigned(16#47#, 8);
  gmul3_9(61) <= to_unsigned(16#42#, 8);
  gmul3_9(62) <= to_unsigned(16#41#, 8);
  gmul3_9(63) <= to_unsigned(16#C0#, 8);
  gmul3_9(64) <= to_unsigned(16#C3#, 8);
  gmul3_9(65) <= to_unsigned(16#C6#, 8);
  gmul3_9(66) <= to_unsigned(16#C5#, 8);
  gmul3_9(67) <= to_unsigned(16#CC#, 8);
  gmul3_9(68) <= to_unsigned(16#CF#, 8);
  gmul3_9(69) <= to_unsigned(16#CA#, 8);
  gmul3_9(70) <= to_unsigned(16#C9#, 8);
  gmul3_9(71) <= to_unsigned(16#D8#, 8);
  gmul3_9(72) <= to_unsigned(16#DB#, 8);
  gmul3_9(73) <= to_unsigned(16#DE#, 8);
  gmul3_9(74) <= to_unsigned(16#DD#, 8);
  gmul3_9(75) <= to_unsigned(16#D4#, 8);
  gmul3_9(76) <= to_unsigned(16#D7#, 8);
  gmul3_9(77) <= to_unsigned(16#D2#, 8);
  gmul3_9(78) <= to_unsigned(16#D1#, 8);
  gmul3_9(79) <= to_unsigned(16#F0#, 8);
  gmul3_9(80) <= to_unsigned(16#F3#, 8);
  gmul3_9(81) <= to_unsigned(16#F6#, 8);
  gmul3_9(82) <= to_unsigned(16#F5#, 8);
  gmul3_9(83) <= to_unsigned(16#FC#, 8);
  gmul3_9(84) <= to_unsigned(16#FF#, 8);
  gmul3_9(85) <= to_unsigned(16#FA#, 8);
  gmul3_9(86) <= to_unsigned(16#F9#, 8);
  gmul3_9(87) <= to_unsigned(16#E8#, 8);
  gmul3_9(88) <= to_unsigned(16#EB#, 8);
  gmul3_9(89) <= to_unsigned(16#EE#, 8);
  gmul3_9(90) <= to_unsigned(16#ED#, 8);
  gmul3_9(91) <= to_unsigned(16#E4#, 8);
  gmul3_9(92) <= to_unsigned(16#E7#, 8);
  gmul3_9(93) <= to_unsigned(16#E2#, 8);
  gmul3_9(94) <= to_unsigned(16#E1#, 8);
  gmul3_9(95) <= to_unsigned(16#A0#, 8);
  gmul3_9(96) <= to_unsigned(16#A3#, 8);
  gmul3_9(97) <= to_unsigned(16#A6#, 8);
  gmul3_9(98) <= to_unsigned(16#A5#, 8);
  gmul3_9(99) <= to_unsigned(16#AC#, 8);
  gmul3_9(100) <= to_unsigned(16#AF#, 8);
  gmul3_9(101) <= to_unsigned(16#AA#, 8);
  gmul3_9(102) <= to_unsigned(16#A9#, 8);
  gmul3_9(103) <= to_unsigned(16#B8#, 8);
  gmul3_9(104) <= to_unsigned(16#BB#, 8);
  gmul3_9(105) <= to_unsigned(16#BE#, 8);
  gmul3_9(106) <= to_unsigned(16#BD#, 8);
  gmul3_9(107) <= to_unsigned(16#B4#, 8);
  gmul3_9(108) <= to_unsigned(16#B7#, 8);
  gmul3_9(109) <= to_unsigned(16#B2#, 8);
  gmul3_9(110) <= to_unsigned(16#B1#, 8);
  gmul3_9(111) <= to_unsigned(16#90#, 8);
  gmul3_9(112) <= to_unsigned(16#93#, 8);
  gmul3_9(113) <= to_unsigned(16#96#, 8);
  gmul3_9(114) <= to_unsigned(16#95#, 8);
  gmul3_9(115) <= to_unsigned(16#9C#, 8);
  gmul3_9(116) <= to_unsigned(16#9F#, 8);
  gmul3_9(117) <= to_unsigned(16#9A#, 8);
  gmul3_9(118) <= to_unsigned(16#99#, 8);
  gmul3_9(119) <= to_unsigned(16#88#, 8);
  gmul3_9(120) <= to_unsigned(16#8B#, 8);
  gmul3_9(121) <= to_unsigned(16#8E#, 8);
  gmul3_9(122) <= to_unsigned(16#8D#, 8);
  gmul3_9(123) <= to_unsigned(16#84#, 8);
  gmul3_9(124) <= to_unsigned(16#87#, 8);
  gmul3_9(125) <= to_unsigned(16#82#, 8);
  gmul3_9(126) <= to_unsigned(16#81#, 8);
  gmul3_9(127) <= to_unsigned(16#9B#, 8);
  gmul3_9(128) <= to_unsigned(16#98#, 8);
  gmul3_9(129) <= to_unsigned(16#9D#, 8);
  gmul3_9(130) <= to_unsigned(16#9E#, 8);
  gmul3_9(131) <= to_unsigned(16#97#, 8);
  gmul3_9(132) <= to_unsigned(16#94#, 8);
  gmul3_9(133) <= to_unsigned(16#91#, 8);
  gmul3_9(134) <= to_unsigned(16#92#, 8);
  gmul3_9(135) <= to_unsigned(16#83#, 8);
  gmul3_9(136) <= to_unsigned(16#80#, 8);
  gmul3_9(137) <= to_unsigned(16#85#, 8);
  gmul3_9(138) <= to_unsigned(16#86#, 8);
  gmul3_9(139) <= to_unsigned(16#8F#, 8);
  gmul3_9(140) <= to_unsigned(16#8C#, 8);
  gmul3_9(141) <= to_unsigned(16#89#, 8);
  gmul3_9(142) <= to_unsigned(16#8A#, 8);
  gmul3_9(143) <= to_unsigned(16#AB#, 8);
  gmul3_9(144) <= to_unsigned(16#A8#, 8);
  gmul3_9(145) <= to_unsigned(16#AD#, 8);
  gmul3_9(146) <= to_unsigned(16#AE#, 8);
  gmul3_9(147) <= to_unsigned(16#A7#, 8);
  gmul3_9(148) <= to_unsigned(16#A4#, 8);
  gmul3_9(149) <= to_unsigned(16#A1#, 8);
  gmul3_9(150) <= to_unsigned(16#A2#, 8);
  gmul3_9(151) <= to_unsigned(16#B3#, 8);
  gmul3_9(152) <= to_unsigned(16#B0#, 8);
  gmul3_9(153) <= to_unsigned(16#B5#, 8);
  gmul3_9(154) <= to_unsigned(16#B6#, 8);
  gmul3_9(155) <= to_unsigned(16#BF#, 8);
  gmul3_9(156) <= to_unsigned(16#BC#, 8);
  gmul3_9(157) <= to_unsigned(16#B9#, 8);
  gmul3_9(158) <= to_unsigned(16#BA#, 8);
  gmul3_9(159) <= to_unsigned(16#FB#, 8);
  gmul3_9(160) <= to_unsigned(16#F8#, 8);
  gmul3_9(161) <= to_unsigned(16#FD#, 8);
  gmul3_9(162) <= to_unsigned(16#FE#, 8);
  gmul3_9(163) <= to_unsigned(16#F7#, 8);
  gmul3_9(164) <= to_unsigned(16#F4#, 8);
  gmul3_9(165) <= to_unsigned(16#F1#, 8);
  gmul3_9(166) <= to_unsigned(16#F2#, 8);
  gmul3_9(167) <= to_unsigned(16#E3#, 8);
  gmul3_9(168) <= to_unsigned(16#E0#, 8);
  gmul3_9(169) <= to_unsigned(16#E5#, 8);
  gmul3_9(170) <= to_unsigned(16#E6#, 8);
  gmul3_9(171) <= to_unsigned(16#EF#, 8);
  gmul3_9(172) <= to_unsigned(16#EC#, 8);
  gmul3_9(173) <= to_unsigned(16#E9#, 8);
  gmul3_9(174) <= to_unsigned(16#EA#, 8);
  gmul3_9(175) <= to_unsigned(16#CB#, 8);
  gmul3_9(176) <= to_unsigned(16#C8#, 8);
  gmul3_9(177) <= to_unsigned(16#CD#, 8);
  gmul3_9(178) <= to_unsigned(16#CE#, 8);
  gmul3_9(179) <= to_unsigned(16#C7#, 8);
  gmul3_9(180) <= to_unsigned(16#C4#, 8);
  gmul3_9(181) <= to_unsigned(16#C1#, 8);
  gmul3_9(182) <= to_unsigned(16#C2#, 8);
  gmul3_9(183) <= to_unsigned(16#D3#, 8);
  gmul3_9(184) <= to_unsigned(16#D0#, 8);
  gmul3_9(185) <= to_unsigned(16#D5#, 8);
  gmul3_9(186) <= to_unsigned(16#D6#, 8);
  gmul3_9(187) <= to_unsigned(16#DF#, 8);
  gmul3_9(188) <= to_unsigned(16#DC#, 8);
  gmul3_9(189) <= to_unsigned(16#D9#, 8);
  gmul3_9(190) <= to_unsigned(16#DA#, 8);
  gmul3_9(191) <= to_unsigned(16#5B#, 8);
  gmul3_9(192) <= to_unsigned(16#58#, 8);
  gmul3_9(193) <= to_unsigned(16#5D#, 8);
  gmul3_9(194) <= to_unsigned(16#5E#, 8);
  gmul3_9(195) <= to_unsigned(16#57#, 8);
  gmul3_9(196) <= to_unsigned(16#54#, 8);
  gmul3_9(197) <= to_unsigned(16#51#, 8);
  gmul3_9(198) <= to_unsigned(16#52#, 8);
  gmul3_9(199) <= to_unsigned(16#43#, 8);
  gmul3_9(200) <= to_unsigned(16#40#, 8);
  gmul3_9(201) <= to_unsigned(16#45#, 8);
  gmul3_9(202) <= to_unsigned(16#46#, 8);
  gmul3_9(203) <= to_unsigned(16#4F#, 8);
  gmul3_9(204) <= to_unsigned(16#4C#, 8);
  gmul3_9(205) <= to_unsigned(16#49#, 8);
  gmul3_9(206) <= to_unsigned(16#4A#, 8);
  gmul3_9(207) <= to_unsigned(16#6B#, 8);
  gmul3_9(208) <= to_unsigned(16#68#, 8);
  gmul3_9(209) <= to_unsigned(16#6D#, 8);
  gmul3_9(210) <= to_unsigned(16#6E#, 8);
  gmul3_9(211) <= to_unsigned(16#67#, 8);
  gmul3_9(212) <= to_unsigned(16#64#, 8);
  gmul3_9(213) <= to_unsigned(16#61#, 8);
  gmul3_9(214) <= to_unsigned(16#62#, 8);
  gmul3_9(215) <= to_unsigned(16#73#, 8);
  gmul3_9(216) <= to_unsigned(16#70#, 8);
  gmul3_9(217) <= to_unsigned(16#75#, 8);
  gmul3_9(218) <= to_unsigned(16#76#, 8);
  gmul3_9(219) <= to_unsigned(16#7F#, 8);
  gmul3_9(220) <= to_unsigned(16#7C#, 8);
  gmul3_9(221) <= to_unsigned(16#79#, 8);
  gmul3_9(222) <= to_unsigned(16#7A#, 8);
  gmul3_9(223) <= to_unsigned(16#3B#, 8);
  gmul3_9(224) <= to_unsigned(16#38#, 8);
  gmul3_9(225) <= to_unsigned(16#3D#, 8);
  gmul3_9(226) <= to_unsigned(16#3E#, 8);
  gmul3_9(227) <= to_unsigned(16#37#, 8);
  gmul3_9(228) <= to_unsigned(16#34#, 8);
  gmul3_9(229) <= to_unsigned(16#31#, 8);
  gmul3_9(230) <= to_unsigned(16#32#, 8);
  gmul3_9(231) <= to_unsigned(16#23#, 8);
  gmul3_9(232) <= to_unsigned(16#20#, 8);
  gmul3_9(233) <= to_unsigned(16#25#, 8);
  gmul3_9(234) <= to_unsigned(16#26#, 8);
  gmul3_9(235) <= to_unsigned(16#2F#, 8);
  gmul3_9(236) <= to_unsigned(16#2C#, 8);
  gmul3_9(237) <= to_unsigned(16#29#, 8);
  gmul3_9(238) <= to_unsigned(16#2A#, 8);
  gmul3_9(239) <= to_unsigned(16#0B#, 8);
  gmul3_9(240) <= to_unsigned(16#08#, 8);
  gmul3_9(241) <= to_unsigned(16#0D#, 8);
  gmul3_9(242) <= to_unsigned(16#0E#, 8);
  gmul3_9(243) <= to_unsigned(16#07#, 8);
  gmul3_9(244) <= to_unsigned(16#04#, 8);
  gmul3_9(245) <= to_unsigned(16#01#, 8);
  gmul3_9(246) <= to_unsigned(16#02#, 8);
  gmul3_9(247) <= to_unsigned(16#13#, 8);
  gmul3_9(248) <= to_unsigned(16#10#, 8);
  gmul3_9(249) <= to_unsigned(16#15#, 8);
  gmul3_9(250) <= to_unsigned(16#16#, 8);
  gmul3_9(251) <= to_unsigned(16#1F#, 8);
  gmul3_9(252) <= to_unsigned(16#1C#, 8);
  gmul3_9(253) <= to_unsigned(16#19#, 8);
  gmul3_9(254) <= to_unsigned(16#1A#, 8);
  gmul3_9(255) <= to_unsigned(16#1A#, 8);

  gmul2_10(0) <= to_unsigned(16#02#, 8);
  gmul2_10(1) <= to_unsigned(16#04#, 8);
  gmul2_10(2) <= to_unsigned(16#06#, 8);
  gmul2_10(3) <= to_unsigned(16#08#, 8);
  gmul2_10(4) <= to_unsigned(16#0A#, 8);
  gmul2_10(5) <= to_unsigned(16#0C#, 8);
  gmul2_10(6) <= to_unsigned(16#0E#, 8);
  gmul2_10(7) <= to_unsigned(16#10#, 8);
  gmul2_10(8) <= to_unsigned(16#12#, 8);
  gmul2_10(9) <= to_unsigned(16#14#, 8);
  gmul2_10(10) <= to_unsigned(16#16#, 8);
  gmul2_10(11) <= to_unsigned(16#18#, 8);
  gmul2_10(12) <= to_unsigned(16#1A#, 8);
  gmul2_10(13) <= to_unsigned(16#1C#, 8);
  gmul2_10(14) <= to_unsigned(16#1E#, 8);
  gmul2_10(15) <= to_unsigned(16#20#, 8);
  gmul2_10(16) <= to_unsigned(16#22#, 8);
  gmul2_10(17) <= to_unsigned(16#24#, 8);
  gmul2_10(18) <= to_unsigned(16#26#, 8);
  gmul2_10(19) <= to_unsigned(16#28#, 8);
  gmul2_10(20) <= to_unsigned(16#2A#, 8);
  gmul2_10(21) <= to_unsigned(16#2C#, 8);
  gmul2_10(22) <= to_unsigned(16#2E#, 8);
  gmul2_10(23) <= to_unsigned(16#30#, 8);
  gmul2_10(24) <= to_unsigned(16#32#, 8);
  gmul2_10(25) <= to_unsigned(16#34#, 8);
  gmul2_10(26) <= to_unsigned(16#36#, 8);
  gmul2_10(27) <= to_unsigned(16#38#, 8);
  gmul2_10(28) <= to_unsigned(16#3A#, 8);
  gmul2_10(29) <= to_unsigned(16#3C#, 8);
  gmul2_10(30) <= to_unsigned(16#3E#, 8);
  gmul2_10(31) <= to_unsigned(16#40#, 8);
  gmul2_10(32) <= to_unsigned(16#42#, 8);
  gmul2_10(33) <= to_unsigned(16#44#, 8);
  gmul2_10(34) <= to_unsigned(16#46#, 8);
  gmul2_10(35) <= to_unsigned(16#48#, 8);
  gmul2_10(36) <= to_unsigned(16#4A#, 8);
  gmul2_10(37) <= to_unsigned(16#4C#, 8);
  gmul2_10(38) <= to_unsigned(16#4E#, 8);
  gmul2_10(39) <= to_unsigned(16#50#, 8);
  gmul2_10(40) <= to_unsigned(16#52#, 8);
  gmul2_10(41) <= to_unsigned(16#54#, 8);
  gmul2_10(42) <= to_unsigned(16#56#, 8);
  gmul2_10(43) <= to_unsigned(16#58#, 8);
  gmul2_10(44) <= to_unsigned(16#5A#, 8);
  gmul2_10(45) <= to_unsigned(16#5C#, 8);
  gmul2_10(46) <= to_unsigned(16#5E#, 8);
  gmul2_10(47) <= to_unsigned(16#60#, 8);
  gmul2_10(48) <= to_unsigned(16#62#, 8);
  gmul2_10(49) <= to_unsigned(16#64#, 8);
  gmul2_10(50) <= to_unsigned(16#66#, 8);
  gmul2_10(51) <= to_unsigned(16#68#, 8);
  gmul2_10(52) <= to_unsigned(16#6A#, 8);
  gmul2_10(53) <= to_unsigned(16#6C#, 8);
  gmul2_10(54) <= to_unsigned(16#6E#, 8);
  gmul2_10(55) <= to_unsigned(16#70#, 8);
  gmul2_10(56) <= to_unsigned(16#72#, 8);
  gmul2_10(57) <= to_unsigned(16#74#, 8);
  gmul2_10(58) <= to_unsigned(16#76#, 8);
  gmul2_10(59) <= to_unsigned(16#78#, 8);
  gmul2_10(60) <= to_unsigned(16#7A#, 8);
  gmul2_10(61) <= to_unsigned(16#7C#, 8);
  gmul2_10(62) <= to_unsigned(16#7E#, 8);
  gmul2_10(63) <= to_unsigned(16#80#, 8);
  gmul2_10(64) <= to_unsigned(16#82#, 8);
  gmul2_10(65) <= to_unsigned(16#84#, 8);
  gmul2_10(66) <= to_unsigned(16#86#, 8);
  gmul2_10(67) <= to_unsigned(16#88#, 8);
  gmul2_10(68) <= to_unsigned(16#8A#, 8);
  gmul2_10(69) <= to_unsigned(16#8C#, 8);
  gmul2_10(70) <= to_unsigned(16#8E#, 8);
  gmul2_10(71) <= to_unsigned(16#90#, 8);
  gmul2_10(72) <= to_unsigned(16#92#, 8);
  gmul2_10(73) <= to_unsigned(16#94#, 8);
  gmul2_10(74) <= to_unsigned(16#96#, 8);
  gmul2_10(75) <= to_unsigned(16#98#, 8);
  gmul2_10(76) <= to_unsigned(16#9A#, 8);
  gmul2_10(77) <= to_unsigned(16#9C#, 8);
  gmul2_10(78) <= to_unsigned(16#9E#, 8);
  gmul2_10(79) <= to_unsigned(16#A0#, 8);
  gmul2_10(80) <= to_unsigned(16#A2#, 8);
  gmul2_10(81) <= to_unsigned(16#A4#, 8);
  gmul2_10(82) <= to_unsigned(16#A6#, 8);
  gmul2_10(83) <= to_unsigned(16#A8#, 8);
  gmul2_10(84) <= to_unsigned(16#AA#, 8);
  gmul2_10(85) <= to_unsigned(16#AC#, 8);
  gmul2_10(86) <= to_unsigned(16#AE#, 8);
  gmul2_10(87) <= to_unsigned(16#B0#, 8);
  gmul2_10(88) <= to_unsigned(16#B2#, 8);
  gmul2_10(89) <= to_unsigned(16#B4#, 8);
  gmul2_10(90) <= to_unsigned(16#B6#, 8);
  gmul2_10(91) <= to_unsigned(16#B8#, 8);
  gmul2_10(92) <= to_unsigned(16#BA#, 8);
  gmul2_10(93) <= to_unsigned(16#BC#, 8);
  gmul2_10(94) <= to_unsigned(16#BE#, 8);
  gmul2_10(95) <= to_unsigned(16#C0#, 8);
  gmul2_10(96) <= to_unsigned(16#C2#, 8);
  gmul2_10(97) <= to_unsigned(16#C4#, 8);
  gmul2_10(98) <= to_unsigned(16#C6#, 8);
  gmul2_10(99) <= to_unsigned(16#C8#, 8);
  gmul2_10(100) <= to_unsigned(16#CA#, 8);
  gmul2_10(101) <= to_unsigned(16#CC#, 8);
  gmul2_10(102) <= to_unsigned(16#CE#, 8);
  gmul2_10(103) <= to_unsigned(16#D0#, 8);
  gmul2_10(104) <= to_unsigned(16#D2#, 8);
  gmul2_10(105) <= to_unsigned(16#D4#, 8);
  gmul2_10(106) <= to_unsigned(16#D6#, 8);
  gmul2_10(107) <= to_unsigned(16#D8#, 8);
  gmul2_10(108) <= to_unsigned(16#DA#, 8);
  gmul2_10(109) <= to_unsigned(16#DC#, 8);
  gmul2_10(110) <= to_unsigned(16#DE#, 8);
  gmul2_10(111) <= to_unsigned(16#E0#, 8);
  gmul2_10(112) <= to_unsigned(16#E2#, 8);
  gmul2_10(113) <= to_unsigned(16#E4#, 8);
  gmul2_10(114) <= to_unsigned(16#E6#, 8);
  gmul2_10(115) <= to_unsigned(16#E8#, 8);
  gmul2_10(116) <= to_unsigned(16#EA#, 8);
  gmul2_10(117) <= to_unsigned(16#EC#, 8);
  gmul2_10(118) <= to_unsigned(16#EE#, 8);
  gmul2_10(119) <= to_unsigned(16#F0#, 8);
  gmul2_10(120) <= to_unsigned(16#F2#, 8);
  gmul2_10(121) <= to_unsigned(16#F4#, 8);
  gmul2_10(122) <= to_unsigned(16#F6#, 8);
  gmul2_10(123) <= to_unsigned(16#F8#, 8);
  gmul2_10(124) <= to_unsigned(16#FA#, 8);
  gmul2_10(125) <= to_unsigned(16#FC#, 8);
  gmul2_10(126) <= to_unsigned(16#FE#, 8);
  gmul2_10(127) <= to_unsigned(16#1B#, 8);
  gmul2_10(128) <= to_unsigned(16#19#, 8);
  gmul2_10(129) <= to_unsigned(16#1F#, 8);
  gmul2_10(130) <= to_unsigned(16#1D#, 8);
  gmul2_10(131) <= to_unsigned(16#13#, 8);
  gmul2_10(132) <= to_unsigned(16#11#, 8);
  gmul2_10(133) <= to_unsigned(16#17#, 8);
  gmul2_10(134) <= to_unsigned(16#15#, 8);
  gmul2_10(135) <= to_unsigned(16#0B#, 8);
  gmul2_10(136) <= to_unsigned(16#09#, 8);
  gmul2_10(137) <= to_unsigned(16#0F#, 8);
  gmul2_10(138) <= to_unsigned(16#0D#, 8);
  gmul2_10(139) <= to_unsigned(16#03#, 8);
  gmul2_10(140) <= to_unsigned(16#01#, 8);
  gmul2_10(141) <= to_unsigned(16#07#, 8);
  gmul2_10(142) <= to_unsigned(16#05#, 8);
  gmul2_10(143) <= to_unsigned(16#3B#, 8);
  gmul2_10(144) <= to_unsigned(16#39#, 8);
  gmul2_10(145) <= to_unsigned(16#3F#, 8);
  gmul2_10(146) <= to_unsigned(16#3D#, 8);
  gmul2_10(147) <= to_unsigned(16#33#, 8);
  gmul2_10(148) <= to_unsigned(16#31#, 8);
  gmul2_10(149) <= to_unsigned(16#37#, 8);
  gmul2_10(150) <= to_unsigned(16#35#, 8);
  gmul2_10(151) <= to_unsigned(16#2B#, 8);
  gmul2_10(152) <= to_unsigned(16#29#, 8);
  gmul2_10(153) <= to_unsigned(16#2F#, 8);
  gmul2_10(154) <= to_unsigned(16#2D#, 8);
  gmul2_10(155) <= to_unsigned(16#23#, 8);
  gmul2_10(156) <= to_unsigned(16#21#, 8);
  gmul2_10(157) <= to_unsigned(16#27#, 8);
  gmul2_10(158) <= to_unsigned(16#25#, 8);
  gmul2_10(159) <= to_unsigned(16#5B#, 8);
  gmul2_10(160) <= to_unsigned(16#59#, 8);
  gmul2_10(161) <= to_unsigned(16#5F#, 8);
  gmul2_10(162) <= to_unsigned(16#5D#, 8);
  gmul2_10(163) <= to_unsigned(16#53#, 8);
  gmul2_10(164) <= to_unsigned(16#51#, 8);
  gmul2_10(165) <= to_unsigned(16#57#, 8);
  gmul2_10(166) <= to_unsigned(16#55#, 8);
  gmul2_10(167) <= to_unsigned(16#4B#, 8);
  gmul2_10(168) <= to_unsigned(16#49#, 8);
  gmul2_10(169) <= to_unsigned(16#4F#, 8);
  gmul2_10(170) <= to_unsigned(16#4D#, 8);
  gmul2_10(171) <= to_unsigned(16#43#, 8);
  gmul2_10(172) <= to_unsigned(16#41#, 8);
  gmul2_10(173) <= to_unsigned(16#47#, 8);
  gmul2_10(174) <= to_unsigned(16#45#, 8);
  gmul2_10(175) <= to_unsigned(16#7B#, 8);
  gmul2_10(176) <= to_unsigned(16#79#, 8);
  gmul2_10(177) <= to_unsigned(16#7F#, 8);
  gmul2_10(178) <= to_unsigned(16#7D#, 8);
  gmul2_10(179) <= to_unsigned(16#73#, 8);
  gmul2_10(180) <= to_unsigned(16#71#, 8);
  gmul2_10(181) <= to_unsigned(16#77#, 8);
  gmul2_10(182) <= to_unsigned(16#75#, 8);
  gmul2_10(183) <= to_unsigned(16#6B#, 8);
  gmul2_10(184) <= to_unsigned(16#69#, 8);
  gmul2_10(185) <= to_unsigned(16#6F#, 8);
  gmul2_10(186) <= to_unsigned(16#6D#, 8);
  gmul2_10(187) <= to_unsigned(16#63#, 8);
  gmul2_10(188) <= to_unsigned(16#61#, 8);
  gmul2_10(189) <= to_unsigned(16#67#, 8);
  gmul2_10(190) <= to_unsigned(16#65#, 8);
  gmul2_10(191) <= to_unsigned(16#9B#, 8);
  gmul2_10(192) <= to_unsigned(16#99#, 8);
  gmul2_10(193) <= to_unsigned(16#9F#, 8);
  gmul2_10(194) <= to_unsigned(16#9D#, 8);
  gmul2_10(195) <= to_unsigned(16#93#, 8);
  gmul2_10(196) <= to_unsigned(16#91#, 8);
  gmul2_10(197) <= to_unsigned(16#97#, 8);
  gmul2_10(198) <= to_unsigned(16#95#, 8);
  gmul2_10(199) <= to_unsigned(16#8B#, 8);
  gmul2_10(200) <= to_unsigned(16#89#, 8);
  gmul2_10(201) <= to_unsigned(16#8F#, 8);
  gmul2_10(202) <= to_unsigned(16#8D#, 8);
  gmul2_10(203) <= to_unsigned(16#83#, 8);
  gmul2_10(204) <= to_unsigned(16#81#, 8);
  gmul2_10(205) <= to_unsigned(16#87#, 8);
  gmul2_10(206) <= to_unsigned(16#85#, 8);
  gmul2_10(207) <= to_unsigned(16#BB#, 8);
  gmul2_10(208) <= to_unsigned(16#B9#, 8);
  gmul2_10(209) <= to_unsigned(16#BF#, 8);
  gmul2_10(210) <= to_unsigned(16#BD#, 8);
  gmul2_10(211) <= to_unsigned(16#B3#, 8);
  gmul2_10(212) <= to_unsigned(16#B1#, 8);
  gmul2_10(213) <= to_unsigned(16#B7#, 8);
  gmul2_10(214) <= to_unsigned(16#B5#, 8);
  gmul2_10(215) <= to_unsigned(16#AB#, 8);
  gmul2_10(216) <= to_unsigned(16#A9#, 8);
  gmul2_10(217) <= to_unsigned(16#AF#, 8);
  gmul2_10(218) <= to_unsigned(16#AD#, 8);
  gmul2_10(219) <= to_unsigned(16#A3#, 8);
  gmul2_10(220) <= to_unsigned(16#A1#, 8);
  gmul2_10(221) <= to_unsigned(16#A7#, 8);
  gmul2_10(222) <= to_unsigned(16#A5#, 8);
  gmul2_10(223) <= to_unsigned(16#DB#, 8);
  gmul2_10(224) <= to_unsigned(16#D9#, 8);
  gmul2_10(225) <= to_unsigned(16#DF#, 8);
  gmul2_10(226) <= to_unsigned(16#DD#, 8);
  gmul2_10(227) <= to_unsigned(16#D3#, 8);
  gmul2_10(228) <= to_unsigned(16#D1#, 8);
  gmul2_10(229) <= to_unsigned(16#D7#, 8);
  gmul2_10(230) <= to_unsigned(16#D5#, 8);
  gmul2_10(231) <= to_unsigned(16#CB#, 8);
  gmul2_10(232) <= to_unsigned(16#C9#, 8);
  gmul2_10(233) <= to_unsigned(16#CF#, 8);
  gmul2_10(234) <= to_unsigned(16#CD#, 8);
  gmul2_10(235) <= to_unsigned(16#C3#, 8);
  gmul2_10(236) <= to_unsigned(16#C1#, 8);
  gmul2_10(237) <= to_unsigned(16#C7#, 8);
  gmul2_10(238) <= to_unsigned(16#C5#, 8);
  gmul2_10(239) <= to_unsigned(16#FB#, 8);
  gmul2_10(240) <= to_unsigned(16#F9#, 8);
  gmul2_10(241) <= to_unsigned(16#FF#, 8);
  gmul2_10(242) <= to_unsigned(16#FD#, 8);
  gmul2_10(243) <= to_unsigned(16#F3#, 8);
  gmul2_10(244) <= to_unsigned(16#F1#, 8);
  gmul2_10(245) <= to_unsigned(16#F7#, 8);
  gmul2_10(246) <= to_unsigned(16#F5#, 8);
  gmul2_10(247) <= to_unsigned(16#EB#, 8);
  gmul2_10(248) <= to_unsigned(16#E9#, 8);
  gmul2_10(249) <= to_unsigned(16#EF#, 8);
  gmul2_10(250) <= to_unsigned(16#ED#, 8);
  gmul2_10(251) <= to_unsigned(16#E3#, 8);
  gmul2_10(252) <= to_unsigned(16#E1#, 8);
  gmul2_10(253) <= to_unsigned(16#E7#, 8);
  gmul2_10(254) <= to_unsigned(16#E5#, 8);
  gmul2_10(255) <= to_unsigned(16#E5#, 8);

  gmul3_10(0) <= to_unsigned(16#03#, 8);
  gmul3_10(1) <= to_unsigned(16#06#, 8);
  gmul3_10(2) <= to_unsigned(16#05#, 8);
  gmul3_10(3) <= to_unsigned(16#0C#, 8);
  gmul3_10(4) <= to_unsigned(16#0F#, 8);
  gmul3_10(5) <= to_unsigned(16#0A#, 8);
  gmul3_10(6) <= to_unsigned(16#09#, 8);
  gmul3_10(7) <= to_unsigned(16#18#, 8);
  gmul3_10(8) <= to_unsigned(16#1B#, 8);
  gmul3_10(9) <= to_unsigned(16#1E#, 8);
  gmul3_10(10) <= to_unsigned(16#1D#, 8);
  gmul3_10(11) <= to_unsigned(16#14#, 8);
  gmul3_10(12) <= to_unsigned(16#17#, 8);
  gmul3_10(13) <= to_unsigned(16#12#, 8);
  gmul3_10(14) <= to_unsigned(16#11#, 8);
  gmul3_10(15) <= to_unsigned(16#30#, 8);
  gmul3_10(16) <= to_unsigned(16#33#, 8);
  gmul3_10(17) <= to_unsigned(16#36#, 8);
  gmul3_10(18) <= to_unsigned(16#35#, 8);
  gmul3_10(19) <= to_unsigned(16#3C#, 8);
  gmul3_10(20) <= to_unsigned(16#3F#, 8);
  gmul3_10(21) <= to_unsigned(16#3A#, 8);
  gmul3_10(22) <= to_unsigned(16#39#, 8);
  gmul3_10(23) <= to_unsigned(16#28#, 8);
  gmul3_10(24) <= to_unsigned(16#2B#, 8);
  gmul3_10(25) <= to_unsigned(16#2E#, 8);
  gmul3_10(26) <= to_unsigned(16#2D#, 8);
  gmul3_10(27) <= to_unsigned(16#24#, 8);
  gmul3_10(28) <= to_unsigned(16#27#, 8);
  gmul3_10(29) <= to_unsigned(16#22#, 8);
  gmul3_10(30) <= to_unsigned(16#21#, 8);
  gmul3_10(31) <= to_unsigned(16#60#, 8);
  gmul3_10(32) <= to_unsigned(16#63#, 8);
  gmul3_10(33) <= to_unsigned(16#66#, 8);
  gmul3_10(34) <= to_unsigned(16#65#, 8);
  gmul3_10(35) <= to_unsigned(16#6C#, 8);
  gmul3_10(36) <= to_unsigned(16#6F#, 8);
  gmul3_10(37) <= to_unsigned(16#6A#, 8);
  gmul3_10(38) <= to_unsigned(16#69#, 8);
  gmul3_10(39) <= to_unsigned(16#78#, 8);
  gmul3_10(40) <= to_unsigned(16#7B#, 8);
  gmul3_10(41) <= to_unsigned(16#7E#, 8);
  gmul3_10(42) <= to_unsigned(16#7D#, 8);
  gmul3_10(43) <= to_unsigned(16#74#, 8);
  gmul3_10(44) <= to_unsigned(16#77#, 8);
  gmul3_10(45) <= to_unsigned(16#72#, 8);
  gmul3_10(46) <= to_unsigned(16#71#, 8);
  gmul3_10(47) <= to_unsigned(16#50#, 8);
  gmul3_10(48) <= to_unsigned(16#53#, 8);
  gmul3_10(49) <= to_unsigned(16#56#, 8);
  gmul3_10(50) <= to_unsigned(16#55#, 8);
  gmul3_10(51) <= to_unsigned(16#5C#, 8);
  gmul3_10(52) <= to_unsigned(16#5F#, 8);
  gmul3_10(53) <= to_unsigned(16#5A#, 8);
  gmul3_10(54) <= to_unsigned(16#59#, 8);
  gmul3_10(55) <= to_unsigned(16#48#, 8);
  gmul3_10(56) <= to_unsigned(16#4B#, 8);
  gmul3_10(57) <= to_unsigned(16#4E#, 8);
  gmul3_10(58) <= to_unsigned(16#4D#, 8);
  gmul3_10(59) <= to_unsigned(16#44#, 8);
  gmul3_10(60) <= to_unsigned(16#47#, 8);
  gmul3_10(61) <= to_unsigned(16#42#, 8);
  gmul3_10(62) <= to_unsigned(16#41#, 8);
  gmul3_10(63) <= to_unsigned(16#C0#, 8);
  gmul3_10(64) <= to_unsigned(16#C3#, 8);
  gmul3_10(65) <= to_unsigned(16#C6#, 8);
  gmul3_10(66) <= to_unsigned(16#C5#, 8);
  gmul3_10(67) <= to_unsigned(16#CC#, 8);
  gmul3_10(68) <= to_unsigned(16#CF#, 8);
  gmul3_10(69) <= to_unsigned(16#CA#, 8);
  gmul3_10(70) <= to_unsigned(16#C9#, 8);
  gmul3_10(71) <= to_unsigned(16#D8#, 8);
  gmul3_10(72) <= to_unsigned(16#DB#, 8);
  gmul3_10(73) <= to_unsigned(16#DE#, 8);
  gmul3_10(74) <= to_unsigned(16#DD#, 8);
  gmul3_10(75) <= to_unsigned(16#D4#, 8);
  gmul3_10(76) <= to_unsigned(16#D7#, 8);
  gmul3_10(77) <= to_unsigned(16#D2#, 8);
  gmul3_10(78) <= to_unsigned(16#D1#, 8);
  gmul3_10(79) <= to_unsigned(16#F0#, 8);
  gmul3_10(80) <= to_unsigned(16#F3#, 8);
  gmul3_10(81) <= to_unsigned(16#F6#, 8);
  gmul3_10(82) <= to_unsigned(16#F5#, 8);
  gmul3_10(83) <= to_unsigned(16#FC#, 8);
  gmul3_10(84) <= to_unsigned(16#FF#, 8);
  gmul3_10(85) <= to_unsigned(16#FA#, 8);
  gmul3_10(86) <= to_unsigned(16#F9#, 8);
  gmul3_10(87) <= to_unsigned(16#E8#, 8);
  gmul3_10(88) <= to_unsigned(16#EB#, 8);
  gmul3_10(89) <= to_unsigned(16#EE#, 8);
  gmul3_10(90) <= to_unsigned(16#ED#, 8);
  gmul3_10(91) <= to_unsigned(16#E4#, 8);
  gmul3_10(92) <= to_unsigned(16#E7#, 8);
  gmul3_10(93) <= to_unsigned(16#E2#, 8);
  gmul3_10(94) <= to_unsigned(16#E1#, 8);
  gmul3_10(95) <= to_unsigned(16#A0#, 8);
  gmul3_10(96) <= to_unsigned(16#A3#, 8);
  gmul3_10(97) <= to_unsigned(16#A6#, 8);
  gmul3_10(98) <= to_unsigned(16#A5#, 8);
  gmul3_10(99) <= to_unsigned(16#AC#, 8);
  gmul3_10(100) <= to_unsigned(16#AF#, 8);
  gmul3_10(101) <= to_unsigned(16#AA#, 8);
  gmul3_10(102) <= to_unsigned(16#A9#, 8);
  gmul3_10(103) <= to_unsigned(16#B8#, 8);
  gmul3_10(104) <= to_unsigned(16#BB#, 8);
  gmul3_10(105) <= to_unsigned(16#BE#, 8);
  gmul3_10(106) <= to_unsigned(16#BD#, 8);
  gmul3_10(107) <= to_unsigned(16#B4#, 8);
  gmul3_10(108) <= to_unsigned(16#B7#, 8);
  gmul3_10(109) <= to_unsigned(16#B2#, 8);
  gmul3_10(110) <= to_unsigned(16#B1#, 8);
  gmul3_10(111) <= to_unsigned(16#90#, 8);
  gmul3_10(112) <= to_unsigned(16#93#, 8);
  gmul3_10(113) <= to_unsigned(16#96#, 8);
  gmul3_10(114) <= to_unsigned(16#95#, 8);
  gmul3_10(115) <= to_unsigned(16#9C#, 8);
  gmul3_10(116) <= to_unsigned(16#9F#, 8);
  gmul3_10(117) <= to_unsigned(16#9A#, 8);
  gmul3_10(118) <= to_unsigned(16#99#, 8);
  gmul3_10(119) <= to_unsigned(16#88#, 8);
  gmul3_10(120) <= to_unsigned(16#8B#, 8);
  gmul3_10(121) <= to_unsigned(16#8E#, 8);
  gmul3_10(122) <= to_unsigned(16#8D#, 8);
  gmul3_10(123) <= to_unsigned(16#84#, 8);
  gmul3_10(124) <= to_unsigned(16#87#, 8);
  gmul3_10(125) <= to_unsigned(16#82#, 8);
  gmul3_10(126) <= to_unsigned(16#81#, 8);
  gmul3_10(127) <= to_unsigned(16#9B#, 8);
  gmul3_10(128) <= to_unsigned(16#98#, 8);
  gmul3_10(129) <= to_unsigned(16#9D#, 8);
  gmul3_10(130) <= to_unsigned(16#9E#, 8);
  gmul3_10(131) <= to_unsigned(16#97#, 8);
  gmul3_10(132) <= to_unsigned(16#94#, 8);
  gmul3_10(133) <= to_unsigned(16#91#, 8);
  gmul3_10(134) <= to_unsigned(16#92#, 8);
  gmul3_10(135) <= to_unsigned(16#83#, 8);
  gmul3_10(136) <= to_unsigned(16#80#, 8);
  gmul3_10(137) <= to_unsigned(16#85#, 8);
  gmul3_10(138) <= to_unsigned(16#86#, 8);
  gmul3_10(139) <= to_unsigned(16#8F#, 8);
  gmul3_10(140) <= to_unsigned(16#8C#, 8);
  gmul3_10(141) <= to_unsigned(16#89#, 8);
  gmul3_10(142) <= to_unsigned(16#8A#, 8);
  gmul3_10(143) <= to_unsigned(16#AB#, 8);
  gmul3_10(144) <= to_unsigned(16#A8#, 8);
  gmul3_10(145) <= to_unsigned(16#AD#, 8);
  gmul3_10(146) <= to_unsigned(16#AE#, 8);
  gmul3_10(147) <= to_unsigned(16#A7#, 8);
  gmul3_10(148) <= to_unsigned(16#A4#, 8);
  gmul3_10(149) <= to_unsigned(16#A1#, 8);
  gmul3_10(150) <= to_unsigned(16#A2#, 8);
  gmul3_10(151) <= to_unsigned(16#B3#, 8);
  gmul3_10(152) <= to_unsigned(16#B0#, 8);
  gmul3_10(153) <= to_unsigned(16#B5#, 8);
  gmul3_10(154) <= to_unsigned(16#B6#, 8);
  gmul3_10(155) <= to_unsigned(16#BF#, 8);
  gmul3_10(156) <= to_unsigned(16#BC#, 8);
  gmul3_10(157) <= to_unsigned(16#B9#, 8);
  gmul3_10(158) <= to_unsigned(16#BA#, 8);
  gmul3_10(159) <= to_unsigned(16#FB#, 8);
  gmul3_10(160) <= to_unsigned(16#F8#, 8);
  gmul3_10(161) <= to_unsigned(16#FD#, 8);
  gmul3_10(162) <= to_unsigned(16#FE#, 8);
  gmul3_10(163) <= to_unsigned(16#F7#, 8);
  gmul3_10(164) <= to_unsigned(16#F4#, 8);
  gmul3_10(165) <= to_unsigned(16#F1#, 8);
  gmul3_10(166) <= to_unsigned(16#F2#, 8);
  gmul3_10(167) <= to_unsigned(16#E3#, 8);
  gmul3_10(168) <= to_unsigned(16#E0#, 8);
  gmul3_10(169) <= to_unsigned(16#E5#, 8);
  gmul3_10(170) <= to_unsigned(16#E6#, 8);
  gmul3_10(171) <= to_unsigned(16#EF#, 8);
  gmul3_10(172) <= to_unsigned(16#EC#, 8);
  gmul3_10(173) <= to_unsigned(16#E9#, 8);
  gmul3_10(174) <= to_unsigned(16#EA#, 8);
  gmul3_10(175) <= to_unsigned(16#CB#, 8);
  gmul3_10(176) <= to_unsigned(16#C8#, 8);
  gmul3_10(177) <= to_unsigned(16#CD#, 8);
  gmul3_10(178) <= to_unsigned(16#CE#, 8);
  gmul3_10(179) <= to_unsigned(16#C7#, 8);
  gmul3_10(180) <= to_unsigned(16#C4#, 8);
  gmul3_10(181) <= to_unsigned(16#C1#, 8);
  gmul3_10(182) <= to_unsigned(16#C2#, 8);
  gmul3_10(183) <= to_unsigned(16#D3#, 8);
  gmul3_10(184) <= to_unsigned(16#D0#, 8);
  gmul3_10(185) <= to_unsigned(16#D5#, 8);
  gmul3_10(186) <= to_unsigned(16#D6#, 8);
  gmul3_10(187) <= to_unsigned(16#DF#, 8);
  gmul3_10(188) <= to_unsigned(16#DC#, 8);
  gmul3_10(189) <= to_unsigned(16#D9#, 8);
  gmul3_10(190) <= to_unsigned(16#DA#, 8);
  gmul3_10(191) <= to_unsigned(16#5B#, 8);
  gmul3_10(192) <= to_unsigned(16#58#, 8);
  gmul3_10(193) <= to_unsigned(16#5D#, 8);
  gmul3_10(194) <= to_unsigned(16#5E#, 8);
  gmul3_10(195) <= to_unsigned(16#57#, 8);
  gmul3_10(196) <= to_unsigned(16#54#, 8);
  gmul3_10(197) <= to_unsigned(16#51#, 8);
  gmul3_10(198) <= to_unsigned(16#52#, 8);
  gmul3_10(199) <= to_unsigned(16#43#, 8);
  gmul3_10(200) <= to_unsigned(16#40#, 8);
  gmul3_10(201) <= to_unsigned(16#45#, 8);
  gmul3_10(202) <= to_unsigned(16#46#, 8);
  gmul3_10(203) <= to_unsigned(16#4F#, 8);
  gmul3_10(204) <= to_unsigned(16#4C#, 8);
  gmul3_10(205) <= to_unsigned(16#49#, 8);
  gmul3_10(206) <= to_unsigned(16#4A#, 8);
  gmul3_10(207) <= to_unsigned(16#6B#, 8);
  gmul3_10(208) <= to_unsigned(16#68#, 8);
  gmul3_10(209) <= to_unsigned(16#6D#, 8);
  gmul3_10(210) <= to_unsigned(16#6E#, 8);
  gmul3_10(211) <= to_unsigned(16#67#, 8);
  gmul3_10(212) <= to_unsigned(16#64#, 8);
  gmul3_10(213) <= to_unsigned(16#61#, 8);
  gmul3_10(214) <= to_unsigned(16#62#, 8);
  gmul3_10(215) <= to_unsigned(16#73#, 8);
  gmul3_10(216) <= to_unsigned(16#70#, 8);
  gmul3_10(217) <= to_unsigned(16#75#, 8);
  gmul3_10(218) <= to_unsigned(16#76#, 8);
  gmul3_10(219) <= to_unsigned(16#7F#, 8);
  gmul3_10(220) <= to_unsigned(16#7C#, 8);
  gmul3_10(221) <= to_unsigned(16#79#, 8);
  gmul3_10(222) <= to_unsigned(16#7A#, 8);
  gmul3_10(223) <= to_unsigned(16#3B#, 8);
  gmul3_10(224) <= to_unsigned(16#38#, 8);
  gmul3_10(225) <= to_unsigned(16#3D#, 8);
  gmul3_10(226) <= to_unsigned(16#3E#, 8);
  gmul3_10(227) <= to_unsigned(16#37#, 8);
  gmul3_10(228) <= to_unsigned(16#34#, 8);
  gmul3_10(229) <= to_unsigned(16#31#, 8);
  gmul3_10(230) <= to_unsigned(16#32#, 8);
  gmul3_10(231) <= to_unsigned(16#23#, 8);
  gmul3_10(232) <= to_unsigned(16#20#, 8);
  gmul3_10(233) <= to_unsigned(16#25#, 8);
  gmul3_10(234) <= to_unsigned(16#26#, 8);
  gmul3_10(235) <= to_unsigned(16#2F#, 8);
  gmul3_10(236) <= to_unsigned(16#2C#, 8);
  gmul3_10(237) <= to_unsigned(16#29#, 8);
  gmul3_10(238) <= to_unsigned(16#2A#, 8);
  gmul3_10(239) <= to_unsigned(16#0B#, 8);
  gmul3_10(240) <= to_unsigned(16#08#, 8);
  gmul3_10(241) <= to_unsigned(16#0D#, 8);
  gmul3_10(242) <= to_unsigned(16#0E#, 8);
  gmul3_10(243) <= to_unsigned(16#07#, 8);
  gmul3_10(244) <= to_unsigned(16#04#, 8);
  gmul3_10(245) <= to_unsigned(16#01#, 8);
  gmul3_10(246) <= to_unsigned(16#02#, 8);
  gmul3_10(247) <= to_unsigned(16#13#, 8);
  gmul3_10(248) <= to_unsigned(16#10#, 8);
  gmul3_10(249) <= to_unsigned(16#15#, 8);
  gmul3_10(250) <= to_unsigned(16#16#, 8);
  gmul3_10(251) <= to_unsigned(16#1F#, 8);
  gmul3_10(252) <= to_unsigned(16#1C#, 8);
  gmul3_10(253) <= to_unsigned(16#19#, 8);
  gmul3_10(254) <= to_unsigned(16#1A#, 8);
  gmul3_10(255) <= to_unsigned(16#1A#, 8);

  gmul3_11(0) <= to_unsigned(16#03#, 8);
  gmul3_11(1) <= to_unsigned(16#06#, 8);
  gmul3_11(2) <= to_unsigned(16#05#, 8);
  gmul3_11(3) <= to_unsigned(16#0C#, 8);
  gmul3_11(4) <= to_unsigned(16#0F#, 8);
  gmul3_11(5) <= to_unsigned(16#0A#, 8);
  gmul3_11(6) <= to_unsigned(16#09#, 8);
  gmul3_11(7) <= to_unsigned(16#18#, 8);
  gmul3_11(8) <= to_unsigned(16#1B#, 8);
  gmul3_11(9) <= to_unsigned(16#1E#, 8);
  gmul3_11(10) <= to_unsigned(16#1D#, 8);
  gmul3_11(11) <= to_unsigned(16#14#, 8);
  gmul3_11(12) <= to_unsigned(16#17#, 8);
  gmul3_11(13) <= to_unsigned(16#12#, 8);
  gmul3_11(14) <= to_unsigned(16#11#, 8);
  gmul3_11(15) <= to_unsigned(16#30#, 8);
  gmul3_11(16) <= to_unsigned(16#33#, 8);
  gmul3_11(17) <= to_unsigned(16#36#, 8);
  gmul3_11(18) <= to_unsigned(16#35#, 8);
  gmul3_11(19) <= to_unsigned(16#3C#, 8);
  gmul3_11(20) <= to_unsigned(16#3F#, 8);
  gmul3_11(21) <= to_unsigned(16#3A#, 8);
  gmul3_11(22) <= to_unsigned(16#39#, 8);
  gmul3_11(23) <= to_unsigned(16#28#, 8);
  gmul3_11(24) <= to_unsigned(16#2B#, 8);
  gmul3_11(25) <= to_unsigned(16#2E#, 8);
  gmul3_11(26) <= to_unsigned(16#2D#, 8);
  gmul3_11(27) <= to_unsigned(16#24#, 8);
  gmul3_11(28) <= to_unsigned(16#27#, 8);
  gmul3_11(29) <= to_unsigned(16#22#, 8);
  gmul3_11(30) <= to_unsigned(16#21#, 8);
  gmul3_11(31) <= to_unsigned(16#60#, 8);
  gmul3_11(32) <= to_unsigned(16#63#, 8);
  gmul3_11(33) <= to_unsigned(16#66#, 8);
  gmul3_11(34) <= to_unsigned(16#65#, 8);
  gmul3_11(35) <= to_unsigned(16#6C#, 8);
  gmul3_11(36) <= to_unsigned(16#6F#, 8);
  gmul3_11(37) <= to_unsigned(16#6A#, 8);
  gmul3_11(38) <= to_unsigned(16#69#, 8);
  gmul3_11(39) <= to_unsigned(16#78#, 8);
  gmul3_11(40) <= to_unsigned(16#7B#, 8);
  gmul3_11(41) <= to_unsigned(16#7E#, 8);
  gmul3_11(42) <= to_unsigned(16#7D#, 8);
  gmul3_11(43) <= to_unsigned(16#74#, 8);
  gmul3_11(44) <= to_unsigned(16#77#, 8);
  gmul3_11(45) <= to_unsigned(16#72#, 8);
  gmul3_11(46) <= to_unsigned(16#71#, 8);
  gmul3_11(47) <= to_unsigned(16#50#, 8);
  gmul3_11(48) <= to_unsigned(16#53#, 8);
  gmul3_11(49) <= to_unsigned(16#56#, 8);
  gmul3_11(50) <= to_unsigned(16#55#, 8);
  gmul3_11(51) <= to_unsigned(16#5C#, 8);
  gmul3_11(52) <= to_unsigned(16#5F#, 8);
  gmul3_11(53) <= to_unsigned(16#5A#, 8);
  gmul3_11(54) <= to_unsigned(16#59#, 8);
  gmul3_11(55) <= to_unsigned(16#48#, 8);
  gmul3_11(56) <= to_unsigned(16#4B#, 8);
  gmul3_11(57) <= to_unsigned(16#4E#, 8);
  gmul3_11(58) <= to_unsigned(16#4D#, 8);
  gmul3_11(59) <= to_unsigned(16#44#, 8);
  gmul3_11(60) <= to_unsigned(16#47#, 8);
  gmul3_11(61) <= to_unsigned(16#42#, 8);
  gmul3_11(62) <= to_unsigned(16#41#, 8);
  gmul3_11(63) <= to_unsigned(16#C0#, 8);
  gmul3_11(64) <= to_unsigned(16#C3#, 8);
  gmul3_11(65) <= to_unsigned(16#C6#, 8);
  gmul3_11(66) <= to_unsigned(16#C5#, 8);
  gmul3_11(67) <= to_unsigned(16#CC#, 8);
  gmul3_11(68) <= to_unsigned(16#CF#, 8);
  gmul3_11(69) <= to_unsigned(16#CA#, 8);
  gmul3_11(70) <= to_unsigned(16#C9#, 8);
  gmul3_11(71) <= to_unsigned(16#D8#, 8);
  gmul3_11(72) <= to_unsigned(16#DB#, 8);
  gmul3_11(73) <= to_unsigned(16#DE#, 8);
  gmul3_11(74) <= to_unsigned(16#DD#, 8);
  gmul3_11(75) <= to_unsigned(16#D4#, 8);
  gmul3_11(76) <= to_unsigned(16#D7#, 8);
  gmul3_11(77) <= to_unsigned(16#D2#, 8);
  gmul3_11(78) <= to_unsigned(16#D1#, 8);
  gmul3_11(79) <= to_unsigned(16#F0#, 8);
  gmul3_11(80) <= to_unsigned(16#F3#, 8);
  gmul3_11(81) <= to_unsigned(16#F6#, 8);
  gmul3_11(82) <= to_unsigned(16#F5#, 8);
  gmul3_11(83) <= to_unsigned(16#FC#, 8);
  gmul3_11(84) <= to_unsigned(16#FF#, 8);
  gmul3_11(85) <= to_unsigned(16#FA#, 8);
  gmul3_11(86) <= to_unsigned(16#F9#, 8);
  gmul3_11(87) <= to_unsigned(16#E8#, 8);
  gmul3_11(88) <= to_unsigned(16#EB#, 8);
  gmul3_11(89) <= to_unsigned(16#EE#, 8);
  gmul3_11(90) <= to_unsigned(16#ED#, 8);
  gmul3_11(91) <= to_unsigned(16#E4#, 8);
  gmul3_11(92) <= to_unsigned(16#E7#, 8);
  gmul3_11(93) <= to_unsigned(16#E2#, 8);
  gmul3_11(94) <= to_unsigned(16#E1#, 8);
  gmul3_11(95) <= to_unsigned(16#A0#, 8);
  gmul3_11(96) <= to_unsigned(16#A3#, 8);
  gmul3_11(97) <= to_unsigned(16#A6#, 8);
  gmul3_11(98) <= to_unsigned(16#A5#, 8);
  gmul3_11(99) <= to_unsigned(16#AC#, 8);
  gmul3_11(100) <= to_unsigned(16#AF#, 8);
  gmul3_11(101) <= to_unsigned(16#AA#, 8);
  gmul3_11(102) <= to_unsigned(16#A9#, 8);
  gmul3_11(103) <= to_unsigned(16#B8#, 8);
  gmul3_11(104) <= to_unsigned(16#BB#, 8);
  gmul3_11(105) <= to_unsigned(16#BE#, 8);
  gmul3_11(106) <= to_unsigned(16#BD#, 8);
  gmul3_11(107) <= to_unsigned(16#B4#, 8);
  gmul3_11(108) <= to_unsigned(16#B7#, 8);
  gmul3_11(109) <= to_unsigned(16#B2#, 8);
  gmul3_11(110) <= to_unsigned(16#B1#, 8);
  gmul3_11(111) <= to_unsigned(16#90#, 8);
  gmul3_11(112) <= to_unsigned(16#93#, 8);
  gmul3_11(113) <= to_unsigned(16#96#, 8);
  gmul3_11(114) <= to_unsigned(16#95#, 8);
  gmul3_11(115) <= to_unsigned(16#9C#, 8);
  gmul3_11(116) <= to_unsigned(16#9F#, 8);
  gmul3_11(117) <= to_unsigned(16#9A#, 8);
  gmul3_11(118) <= to_unsigned(16#99#, 8);
  gmul3_11(119) <= to_unsigned(16#88#, 8);
  gmul3_11(120) <= to_unsigned(16#8B#, 8);
  gmul3_11(121) <= to_unsigned(16#8E#, 8);
  gmul3_11(122) <= to_unsigned(16#8D#, 8);
  gmul3_11(123) <= to_unsigned(16#84#, 8);
  gmul3_11(124) <= to_unsigned(16#87#, 8);
  gmul3_11(125) <= to_unsigned(16#82#, 8);
  gmul3_11(126) <= to_unsigned(16#81#, 8);
  gmul3_11(127) <= to_unsigned(16#9B#, 8);
  gmul3_11(128) <= to_unsigned(16#98#, 8);
  gmul3_11(129) <= to_unsigned(16#9D#, 8);
  gmul3_11(130) <= to_unsigned(16#9E#, 8);
  gmul3_11(131) <= to_unsigned(16#97#, 8);
  gmul3_11(132) <= to_unsigned(16#94#, 8);
  gmul3_11(133) <= to_unsigned(16#91#, 8);
  gmul3_11(134) <= to_unsigned(16#92#, 8);
  gmul3_11(135) <= to_unsigned(16#83#, 8);
  gmul3_11(136) <= to_unsigned(16#80#, 8);
  gmul3_11(137) <= to_unsigned(16#85#, 8);
  gmul3_11(138) <= to_unsigned(16#86#, 8);
  gmul3_11(139) <= to_unsigned(16#8F#, 8);
  gmul3_11(140) <= to_unsigned(16#8C#, 8);
  gmul3_11(141) <= to_unsigned(16#89#, 8);
  gmul3_11(142) <= to_unsigned(16#8A#, 8);
  gmul3_11(143) <= to_unsigned(16#AB#, 8);
  gmul3_11(144) <= to_unsigned(16#A8#, 8);
  gmul3_11(145) <= to_unsigned(16#AD#, 8);
  gmul3_11(146) <= to_unsigned(16#AE#, 8);
  gmul3_11(147) <= to_unsigned(16#A7#, 8);
  gmul3_11(148) <= to_unsigned(16#A4#, 8);
  gmul3_11(149) <= to_unsigned(16#A1#, 8);
  gmul3_11(150) <= to_unsigned(16#A2#, 8);
  gmul3_11(151) <= to_unsigned(16#B3#, 8);
  gmul3_11(152) <= to_unsigned(16#B0#, 8);
  gmul3_11(153) <= to_unsigned(16#B5#, 8);
  gmul3_11(154) <= to_unsigned(16#B6#, 8);
  gmul3_11(155) <= to_unsigned(16#BF#, 8);
  gmul3_11(156) <= to_unsigned(16#BC#, 8);
  gmul3_11(157) <= to_unsigned(16#B9#, 8);
  gmul3_11(158) <= to_unsigned(16#BA#, 8);
  gmul3_11(159) <= to_unsigned(16#FB#, 8);
  gmul3_11(160) <= to_unsigned(16#F8#, 8);
  gmul3_11(161) <= to_unsigned(16#FD#, 8);
  gmul3_11(162) <= to_unsigned(16#FE#, 8);
  gmul3_11(163) <= to_unsigned(16#F7#, 8);
  gmul3_11(164) <= to_unsigned(16#F4#, 8);
  gmul3_11(165) <= to_unsigned(16#F1#, 8);
  gmul3_11(166) <= to_unsigned(16#F2#, 8);
  gmul3_11(167) <= to_unsigned(16#E3#, 8);
  gmul3_11(168) <= to_unsigned(16#E0#, 8);
  gmul3_11(169) <= to_unsigned(16#E5#, 8);
  gmul3_11(170) <= to_unsigned(16#E6#, 8);
  gmul3_11(171) <= to_unsigned(16#EF#, 8);
  gmul3_11(172) <= to_unsigned(16#EC#, 8);
  gmul3_11(173) <= to_unsigned(16#E9#, 8);
  gmul3_11(174) <= to_unsigned(16#EA#, 8);
  gmul3_11(175) <= to_unsigned(16#CB#, 8);
  gmul3_11(176) <= to_unsigned(16#C8#, 8);
  gmul3_11(177) <= to_unsigned(16#CD#, 8);
  gmul3_11(178) <= to_unsigned(16#CE#, 8);
  gmul3_11(179) <= to_unsigned(16#C7#, 8);
  gmul3_11(180) <= to_unsigned(16#C4#, 8);
  gmul3_11(181) <= to_unsigned(16#C1#, 8);
  gmul3_11(182) <= to_unsigned(16#C2#, 8);
  gmul3_11(183) <= to_unsigned(16#D3#, 8);
  gmul3_11(184) <= to_unsigned(16#D0#, 8);
  gmul3_11(185) <= to_unsigned(16#D5#, 8);
  gmul3_11(186) <= to_unsigned(16#D6#, 8);
  gmul3_11(187) <= to_unsigned(16#DF#, 8);
  gmul3_11(188) <= to_unsigned(16#DC#, 8);
  gmul3_11(189) <= to_unsigned(16#D9#, 8);
  gmul3_11(190) <= to_unsigned(16#DA#, 8);
  gmul3_11(191) <= to_unsigned(16#5B#, 8);
  gmul3_11(192) <= to_unsigned(16#58#, 8);
  gmul3_11(193) <= to_unsigned(16#5D#, 8);
  gmul3_11(194) <= to_unsigned(16#5E#, 8);
  gmul3_11(195) <= to_unsigned(16#57#, 8);
  gmul3_11(196) <= to_unsigned(16#54#, 8);
  gmul3_11(197) <= to_unsigned(16#51#, 8);
  gmul3_11(198) <= to_unsigned(16#52#, 8);
  gmul3_11(199) <= to_unsigned(16#43#, 8);
  gmul3_11(200) <= to_unsigned(16#40#, 8);
  gmul3_11(201) <= to_unsigned(16#45#, 8);
  gmul3_11(202) <= to_unsigned(16#46#, 8);
  gmul3_11(203) <= to_unsigned(16#4F#, 8);
  gmul3_11(204) <= to_unsigned(16#4C#, 8);
  gmul3_11(205) <= to_unsigned(16#49#, 8);
  gmul3_11(206) <= to_unsigned(16#4A#, 8);
  gmul3_11(207) <= to_unsigned(16#6B#, 8);
  gmul3_11(208) <= to_unsigned(16#68#, 8);
  gmul3_11(209) <= to_unsigned(16#6D#, 8);
  gmul3_11(210) <= to_unsigned(16#6E#, 8);
  gmul3_11(211) <= to_unsigned(16#67#, 8);
  gmul3_11(212) <= to_unsigned(16#64#, 8);
  gmul3_11(213) <= to_unsigned(16#61#, 8);
  gmul3_11(214) <= to_unsigned(16#62#, 8);
  gmul3_11(215) <= to_unsigned(16#73#, 8);
  gmul3_11(216) <= to_unsigned(16#70#, 8);
  gmul3_11(217) <= to_unsigned(16#75#, 8);
  gmul3_11(218) <= to_unsigned(16#76#, 8);
  gmul3_11(219) <= to_unsigned(16#7F#, 8);
  gmul3_11(220) <= to_unsigned(16#7C#, 8);
  gmul3_11(221) <= to_unsigned(16#79#, 8);
  gmul3_11(222) <= to_unsigned(16#7A#, 8);
  gmul3_11(223) <= to_unsigned(16#3B#, 8);
  gmul3_11(224) <= to_unsigned(16#38#, 8);
  gmul3_11(225) <= to_unsigned(16#3D#, 8);
  gmul3_11(226) <= to_unsigned(16#3E#, 8);
  gmul3_11(227) <= to_unsigned(16#37#, 8);
  gmul3_11(228) <= to_unsigned(16#34#, 8);
  gmul3_11(229) <= to_unsigned(16#31#, 8);
  gmul3_11(230) <= to_unsigned(16#32#, 8);
  gmul3_11(231) <= to_unsigned(16#23#, 8);
  gmul3_11(232) <= to_unsigned(16#20#, 8);
  gmul3_11(233) <= to_unsigned(16#25#, 8);
  gmul3_11(234) <= to_unsigned(16#26#, 8);
  gmul3_11(235) <= to_unsigned(16#2F#, 8);
  gmul3_11(236) <= to_unsigned(16#2C#, 8);
  gmul3_11(237) <= to_unsigned(16#29#, 8);
  gmul3_11(238) <= to_unsigned(16#2A#, 8);
  gmul3_11(239) <= to_unsigned(16#0B#, 8);
  gmul3_11(240) <= to_unsigned(16#08#, 8);
  gmul3_11(241) <= to_unsigned(16#0D#, 8);
  gmul3_11(242) <= to_unsigned(16#0E#, 8);
  gmul3_11(243) <= to_unsigned(16#07#, 8);
  gmul3_11(244) <= to_unsigned(16#04#, 8);
  gmul3_11(245) <= to_unsigned(16#01#, 8);
  gmul3_11(246) <= to_unsigned(16#02#, 8);
  gmul3_11(247) <= to_unsigned(16#13#, 8);
  gmul3_11(248) <= to_unsigned(16#10#, 8);
  gmul3_11(249) <= to_unsigned(16#15#, 8);
  gmul3_11(250) <= to_unsigned(16#16#, 8);
  gmul3_11(251) <= to_unsigned(16#1F#, 8);
  gmul3_11(252) <= to_unsigned(16#1C#, 8);
  gmul3_11(253) <= to_unsigned(16#19#, 8);
  gmul3_11(254) <= to_unsigned(16#1A#, 8);
  gmul3_11(255) <= to_unsigned(16#1A#, 8);

  gmul2_11(0) <= to_unsigned(16#02#, 8);
  gmul2_11(1) <= to_unsigned(16#04#, 8);
  gmul2_11(2) <= to_unsigned(16#06#, 8);
  gmul2_11(3) <= to_unsigned(16#08#, 8);
  gmul2_11(4) <= to_unsigned(16#0A#, 8);
  gmul2_11(5) <= to_unsigned(16#0C#, 8);
  gmul2_11(6) <= to_unsigned(16#0E#, 8);
  gmul2_11(7) <= to_unsigned(16#10#, 8);
  gmul2_11(8) <= to_unsigned(16#12#, 8);
  gmul2_11(9) <= to_unsigned(16#14#, 8);
  gmul2_11(10) <= to_unsigned(16#16#, 8);
  gmul2_11(11) <= to_unsigned(16#18#, 8);
  gmul2_11(12) <= to_unsigned(16#1A#, 8);
  gmul2_11(13) <= to_unsigned(16#1C#, 8);
  gmul2_11(14) <= to_unsigned(16#1E#, 8);
  gmul2_11(15) <= to_unsigned(16#20#, 8);
  gmul2_11(16) <= to_unsigned(16#22#, 8);
  gmul2_11(17) <= to_unsigned(16#24#, 8);
  gmul2_11(18) <= to_unsigned(16#26#, 8);
  gmul2_11(19) <= to_unsigned(16#28#, 8);
  gmul2_11(20) <= to_unsigned(16#2A#, 8);
  gmul2_11(21) <= to_unsigned(16#2C#, 8);
  gmul2_11(22) <= to_unsigned(16#2E#, 8);
  gmul2_11(23) <= to_unsigned(16#30#, 8);
  gmul2_11(24) <= to_unsigned(16#32#, 8);
  gmul2_11(25) <= to_unsigned(16#34#, 8);
  gmul2_11(26) <= to_unsigned(16#36#, 8);
  gmul2_11(27) <= to_unsigned(16#38#, 8);
  gmul2_11(28) <= to_unsigned(16#3A#, 8);
  gmul2_11(29) <= to_unsigned(16#3C#, 8);
  gmul2_11(30) <= to_unsigned(16#3E#, 8);
  gmul2_11(31) <= to_unsigned(16#40#, 8);
  gmul2_11(32) <= to_unsigned(16#42#, 8);
  gmul2_11(33) <= to_unsigned(16#44#, 8);
  gmul2_11(34) <= to_unsigned(16#46#, 8);
  gmul2_11(35) <= to_unsigned(16#48#, 8);
  gmul2_11(36) <= to_unsigned(16#4A#, 8);
  gmul2_11(37) <= to_unsigned(16#4C#, 8);
  gmul2_11(38) <= to_unsigned(16#4E#, 8);
  gmul2_11(39) <= to_unsigned(16#50#, 8);
  gmul2_11(40) <= to_unsigned(16#52#, 8);
  gmul2_11(41) <= to_unsigned(16#54#, 8);
  gmul2_11(42) <= to_unsigned(16#56#, 8);
  gmul2_11(43) <= to_unsigned(16#58#, 8);
  gmul2_11(44) <= to_unsigned(16#5A#, 8);
  gmul2_11(45) <= to_unsigned(16#5C#, 8);
  gmul2_11(46) <= to_unsigned(16#5E#, 8);
  gmul2_11(47) <= to_unsigned(16#60#, 8);
  gmul2_11(48) <= to_unsigned(16#62#, 8);
  gmul2_11(49) <= to_unsigned(16#64#, 8);
  gmul2_11(50) <= to_unsigned(16#66#, 8);
  gmul2_11(51) <= to_unsigned(16#68#, 8);
  gmul2_11(52) <= to_unsigned(16#6A#, 8);
  gmul2_11(53) <= to_unsigned(16#6C#, 8);
  gmul2_11(54) <= to_unsigned(16#6E#, 8);
  gmul2_11(55) <= to_unsigned(16#70#, 8);
  gmul2_11(56) <= to_unsigned(16#72#, 8);
  gmul2_11(57) <= to_unsigned(16#74#, 8);
  gmul2_11(58) <= to_unsigned(16#76#, 8);
  gmul2_11(59) <= to_unsigned(16#78#, 8);
  gmul2_11(60) <= to_unsigned(16#7A#, 8);
  gmul2_11(61) <= to_unsigned(16#7C#, 8);
  gmul2_11(62) <= to_unsigned(16#7E#, 8);
  gmul2_11(63) <= to_unsigned(16#80#, 8);
  gmul2_11(64) <= to_unsigned(16#82#, 8);
  gmul2_11(65) <= to_unsigned(16#84#, 8);
  gmul2_11(66) <= to_unsigned(16#86#, 8);
  gmul2_11(67) <= to_unsigned(16#88#, 8);
  gmul2_11(68) <= to_unsigned(16#8A#, 8);
  gmul2_11(69) <= to_unsigned(16#8C#, 8);
  gmul2_11(70) <= to_unsigned(16#8E#, 8);
  gmul2_11(71) <= to_unsigned(16#90#, 8);
  gmul2_11(72) <= to_unsigned(16#92#, 8);
  gmul2_11(73) <= to_unsigned(16#94#, 8);
  gmul2_11(74) <= to_unsigned(16#96#, 8);
  gmul2_11(75) <= to_unsigned(16#98#, 8);
  gmul2_11(76) <= to_unsigned(16#9A#, 8);
  gmul2_11(77) <= to_unsigned(16#9C#, 8);
  gmul2_11(78) <= to_unsigned(16#9E#, 8);
  gmul2_11(79) <= to_unsigned(16#A0#, 8);
  gmul2_11(80) <= to_unsigned(16#A2#, 8);
  gmul2_11(81) <= to_unsigned(16#A4#, 8);
  gmul2_11(82) <= to_unsigned(16#A6#, 8);
  gmul2_11(83) <= to_unsigned(16#A8#, 8);
  gmul2_11(84) <= to_unsigned(16#AA#, 8);
  gmul2_11(85) <= to_unsigned(16#AC#, 8);
  gmul2_11(86) <= to_unsigned(16#AE#, 8);
  gmul2_11(87) <= to_unsigned(16#B0#, 8);
  gmul2_11(88) <= to_unsigned(16#B2#, 8);
  gmul2_11(89) <= to_unsigned(16#B4#, 8);
  gmul2_11(90) <= to_unsigned(16#B6#, 8);
  gmul2_11(91) <= to_unsigned(16#B8#, 8);
  gmul2_11(92) <= to_unsigned(16#BA#, 8);
  gmul2_11(93) <= to_unsigned(16#BC#, 8);
  gmul2_11(94) <= to_unsigned(16#BE#, 8);
  gmul2_11(95) <= to_unsigned(16#C0#, 8);
  gmul2_11(96) <= to_unsigned(16#C2#, 8);
  gmul2_11(97) <= to_unsigned(16#C4#, 8);
  gmul2_11(98) <= to_unsigned(16#C6#, 8);
  gmul2_11(99) <= to_unsigned(16#C8#, 8);
  gmul2_11(100) <= to_unsigned(16#CA#, 8);
  gmul2_11(101) <= to_unsigned(16#CC#, 8);
  gmul2_11(102) <= to_unsigned(16#CE#, 8);
  gmul2_11(103) <= to_unsigned(16#D0#, 8);
  gmul2_11(104) <= to_unsigned(16#D2#, 8);
  gmul2_11(105) <= to_unsigned(16#D4#, 8);
  gmul2_11(106) <= to_unsigned(16#D6#, 8);
  gmul2_11(107) <= to_unsigned(16#D8#, 8);
  gmul2_11(108) <= to_unsigned(16#DA#, 8);
  gmul2_11(109) <= to_unsigned(16#DC#, 8);
  gmul2_11(110) <= to_unsigned(16#DE#, 8);
  gmul2_11(111) <= to_unsigned(16#E0#, 8);
  gmul2_11(112) <= to_unsigned(16#E2#, 8);
  gmul2_11(113) <= to_unsigned(16#E4#, 8);
  gmul2_11(114) <= to_unsigned(16#E6#, 8);
  gmul2_11(115) <= to_unsigned(16#E8#, 8);
  gmul2_11(116) <= to_unsigned(16#EA#, 8);
  gmul2_11(117) <= to_unsigned(16#EC#, 8);
  gmul2_11(118) <= to_unsigned(16#EE#, 8);
  gmul2_11(119) <= to_unsigned(16#F0#, 8);
  gmul2_11(120) <= to_unsigned(16#F2#, 8);
  gmul2_11(121) <= to_unsigned(16#F4#, 8);
  gmul2_11(122) <= to_unsigned(16#F6#, 8);
  gmul2_11(123) <= to_unsigned(16#F8#, 8);
  gmul2_11(124) <= to_unsigned(16#FA#, 8);
  gmul2_11(125) <= to_unsigned(16#FC#, 8);
  gmul2_11(126) <= to_unsigned(16#FE#, 8);
  gmul2_11(127) <= to_unsigned(16#1B#, 8);
  gmul2_11(128) <= to_unsigned(16#19#, 8);
  gmul2_11(129) <= to_unsigned(16#1F#, 8);
  gmul2_11(130) <= to_unsigned(16#1D#, 8);
  gmul2_11(131) <= to_unsigned(16#13#, 8);
  gmul2_11(132) <= to_unsigned(16#11#, 8);
  gmul2_11(133) <= to_unsigned(16#17#, 8);
  gmul2_11(134) <= to_unsigned(16#15#, 8);
  gmul2_11(135) <= to_unsigned(16#0B#, 8);
  gmul2_11(136) <= to_unsigned(16#09#, 8);
  gmul2_11(137) <= to_unsigned(16#0F#, 8);
  gmul2_11(138) <= to_unsigned(16#0D#, 8);
  gmul2_11(139) <= to_unsigned(16#03#, 8);
  gmul2_11(140) <= to_unsigned(16#01#, 8);
  gmul2_11(141) <= to_unsigned(16#07#, 8);
  gmul2_11(142) <= to_unsigned(16#05#, 8);
  gmul2_11(143) <= to_unsigned(16#3B#, 8);
  gmul2_11(144) <= to_unsigned(16#39#, 8);
  gmul2_11(145) <= to_unsigned(16#3F#, 8);
  gmul2_11(146) <= to_unsigned(16#3D#, 8);
  gmul2_11(147) <= to_unsigned(16#33#, 8);
  gmul2_11(148) <= to_unsigned(16#31#, 8);
  gmul2_11(149) <= to_unsigned(16#37#, 8);
  gmul2_11(150) <= to_unsigned(16#35#, 8);
  gmul2_11(151) <= to_unsigned(16#2B#, 8);
  gmul2_11(152) <= to_unsigned(16#29#, 8);
  gmul2_11(153) <= to_unsigned(16#2F#, 8);
  gmul2_11(154) <= to_unsigned(16#2D#, 8);
  gmul2_11(155) <= to_unsigned(16#23#, 8);
  gmul2_11(156) <= to_unsigned(16#21#, 8);
  gmul2_11(157) <= to_unsigned(16#27#, 8);
  gmul2_11(158) <= to_unsigned(16#25#, 8);
  gmul2_11(159) <= to_unsigned(16#5B#, 8);
  gmul2_11(160) <= to_unsigned(16#59#, 8);
  gmul2_11(161) <= to_unsigned(16#5F#, 8);
  gmul2_11(162) <= to_unsigned(16#5D#, 8);
  gmul2_11(163) <= to_unsigned(16#53#, 8);
  gmul2_11(164) <= to_unsigned(16#51#, 8);
  gmul2_11(165) <= to_unsigned(16#57#, 8);
  gmul2_11(166) <= to_unsigned(16#55#, 8);
  gmul2_11(167) <= to_unsigned(16#4B#, 8);
  gmul2_11(168) <= to_unsigned(16#49#, 8);
  gmul2_11(169) <= to_unsigned(16#4F#, 8);
  gmul2_11(170) <= to_unsigned(16#4D#, 8);
  gmul2_11(171) <= to_unsigned(16#43#, 8);
  gmul2_11(172) <= to_unsigned(16#41#, 8);
  gmul2_11(173) <= to_unsigned(16#47#, 8);
  gmul2_11(174) <= to_unsigned(16#45#, 8);
  gmul2_11(175) <= to_unsigned(16#7B#, 8);
  gmul2_11(176) <= to_unsigned(16#79#, 8);
  gmul2_11(177) <= to_unsigned(16#7F#, 8);
  gmul2_11(178) <= to_unsigned(16#7D#, 8);
  gmul2_11(179) <= to_unsigned(16#73#, 8);
  gmul2_11(180) <= to_unsigned(16#71#, 8);
  gmul2_11(181) <= to_unsigned(16#77#, 8);
  gmul2_11(182) <= to_unsigned(16#75#, 8);
  gmul2_11(183) <= to_unsigned(16#6B#, 8);
  gmul2_11(184) <= to_unsigned(16#69#, 8);
  gmul2_11(185) <= to_unsigned(16#6F#, 8);
  gmul2_11(186) <= to_unsigned(16#6D#, 8);
  gmul2_11(187) <= to_unsigned(16#63#, 8);
  gmul2_11(188) <= to_unsigned(16#61#, 8);
  gmul2_11(189) <= to_unsigned(16#67#, 8);
  gmul2_11(190) <= to_unsigned(16#65#, 8);
  gmul2_11(191) <= to_unsigned(16#9B#, 8);
  gmul2_11(192) <= to_unsigned(16#99#, 8);
  gmul2_11(193) <= to_unsigned(16#9F#, 8);
  gmul2_11(194) <= to_unsigned(16#9D#, 8);
  gmul2_11(195) <= to_unsigned(16#93#, 8);
  gmul2_11(196) <= to_unsigned(16#91#, 8);
  gmul2_11(197) <= to_unsigned(16#97#, 8);
  gmul2_11(198) <= to_unsigned(16#95#, 8);
  gmul2_11(199) <= to_unsigned(16#8B#, 8);
  gmul2_11(200) <= to_unsigned(16#89#, 8);
  gmul2_11(201) <= to_unsigned(16#8F#, 8);
  gmul2_11(202) <= to_unsigned(16#8D#, 8);
  gmul2_11(203) <= to_unsigned(16#83#, 8);
  gmul2_11(204) <= to_unsigned(16#81#, 8);
  gmul2_11(205) <= to_unsigned(16#87#, 8);
  gmul2_11(206) <= to_unsigned(16#85#, 8);
  gmul2_11(207) <= to_unsigned(16#BB#, 8);
  gmul2_11(208) <= to_unsigned(16#B9#, 8);
  gmul2_11(209) <= to_unsigned(16#BF#, 8);
  gmul2_11(210) <= to_unsigned(16#BD#, 8);
  gmul2_11(211) <= to_unsigned(16#B3#, 8);
  gmul2_11(212) <= to_unsigned(16#B1#, 8);
  gmul2_11(213) <= to_unsigned(16#B7#, 8);
  gmul2_11(214) <= to_unsigned(16#B5#, 8);
  gmul2_11(215) <= to_unsigned(16#AB#, 8);
  gmul2_11(216) <= to_unsigned(16#A9#, 8);
  gmul2_11(217) <= to_unsigned(16#AF#, 8);
  gmul2_11(218) <= to_unsigned(16#AD#, 8);
  gmul2_11(219) <= to_unsigned(16#A3#, 8);
  gmul2_11(220) <= to_unsigned(16#A1#, 8);
  gmul2_11(221) <= to_unsigned(16#A7#, 8);
  gmul2_11(222) <= to_unsigned(16#A5#, 8);
  gmul2_11(223) <= to_unsigned(16#DB#, 8);
  gmul2_11(224) <= to_unsigned(16#D9#, 8);
  gmul2_11(225) <= to_unsigned(16#DF#, 8);
  gmul2_11(226) <= to_unsigned(16#DD#, 8);
  gmul2_11(227) <= to_unsigned(16#D3#, 8);
  gmul2_11(228) <= to_unsigned(16#D1#, 8);
  gmul2_11(229) <= to_unsigned(16#D7#, 8);
  gmul2_11(230) <= to_unsigned(16#D5#, 8);
  gmul2_11(231) <= to_unsigned(16#CB#, 8);
  gmul2_11(232) <= to_unsigned(16#C9#, 8);
  gmul2_11(233) <= to_unsigned(16#CF#, 8);
  gmul2_11(234) <= to_unsigned(16#CD#, 8);
  gmul2_11(235) <= to_unsigned(16#C3#, 8);
  gmul2_11(236) <= to_unsigned(16#C1#, 8);
  gmul2_11(237) <= to_unsigned(16#C7#, 8);
  gmul2_11(238) <= to_unsigned(16#C5#, 8);
  gmul2_11(239) <= to_unsigned(16#FB#, 8);
  gmul2_11(240) <= to_unsigned(16#F9#, 8);
  gmul2_11(241) <= to_unsigned(16#FF#, 8);
  gmul2_11(242) <= to_unsigned(16#FD#, 8);
  gmul2_11(243) <= to_unsigned(16#F3#, 8);
  gmul2_11(244) <= to_unsigned(16#F1#, 8);
  gmul2_11(245) <= to_unsigned(16#F7#, 8);
  gmul2_11(246) <= to_unsigned(16#F5#, 8);
  gmul2_11(247) <= to_unsigned(16#EB#, 8);
  gmul2_11(248) <= to_unsigned(16#E9#, 8);
  gmul2_11(249) <= to_unsigned(16#EF#, 8);
  gmul2_11(250) <= to_unsigned(16#ED#, 8);
  gmul2_11(251) <= to_unsigned(16#E3#, 8);
  gmul2_11(252) <= to_unsigned(16#E1#, 8);
  gmul2_11(253) <= to_unsigned(16#E7#, 8);
  gmul2_11(254) <= to_unsigned(16#E5#, 8);
  gmul2_11(255) <= to_unsigned(16#E5#, 8);

  gmul2_12(0) <= to_unsigned(16#02#, 8);
  gmul2_12(1) <= to_unsigned(16#04#, 8);
  gmul2_12(2) <= to_unsigned(16#06#, 8);
  gmul2_12(3) <= to_unsigned(16#08#, 8);
  gmul2_12(4) <= to_unsigned(16#0A#, 8);
  gmul2_12(5) <= to_unsigned(16#0C#, 8);
  gmul2_12(6) <= to_unsigned(16#0E#, 8);
  gmul2_12(7) <= to_unsigned(16#10#, 8);
  gmul2_12(8) <= to_unsigned(16#12#, 8);
  gmul2_12(9) <= to_unsigned(16#14#, 8);
  gmul2_12(10) <= to_unsigned(16#16#, 8);
  gmul2_12(11) <= to_unsigned(16#18#, 8);
  gmul2_12(12) <= to_unsigned(16#1A#, 8);
  gmul2_12(13) <= to_unsigned(16#1C#, 8);
  gmul2_12(14) <= to_unsigned(16#1E#, 8);
  gmul2_12(15) <= to_unsigned(16#20#, 8);
  gmul2_12(16) <= to_unsigned(16#22#, 8);
  gmul2_12(17) <= to_unsigned(16#24#, 8);
  gmul2_12(18) <= to_unsigned(16#26#, 8);
  gmul2_12(19) <= to_unsigned(16#28#, 8);
  gmul2_12(20) <= to_unsigned(16#2A#, 8);
  gmul2_12(21) <= to_unsigned(16#2C#, 8);
  gmul2_12(22) <= to_unsigned(16#2E#, 8);
  gmul2_12(23) <= to_unsigned(16#30#, 8);
  gmul2_12(24) <= to_unsigned(16#32#, 8);
  gmul2_12(25) <= to_unsigned(16#34#, 8);
  gmul2_12(26) <= to_unsigned(16#36#, 8);
  gmul2_12(27) <= to_unsigned(16#38#, 8);
  gmul2_12(28) <= to_unsigned(16#3A#, 8);
  gmul2_12(29) <= to_unsigned(16#3C#, 8);
  gmul2_12(30) <= to_unsigned(16#3E#, 8);
  gmul2_12(31) <= to_unsigned(16#40#, 8);
  gmul2_12(32) <= to_unsigned(16#42#, 8);
  gmul2_12(33) <= to_unsigned(16#44#, 8);
  gmul2_12(34) <= to_unsigned(16#46#, 8);
  gmul2_12(35) <= to_unsigned(16#48#, 8);
  gmul2_12(36) <= to_unsigned(16#4A#, 8);
  gmul2_12(37) <= to_unsigned(16#4C#, 8);
  gmul2_12(38) <= to_unsigned(16#4E#, 8);
  gmul2_12(39) <= to_unsigned(16#50#, 8);
  gmul2_12(40) <= to_unsigned(16#52#, 8);
  gmul2_12(41) <= to_unsigned(16#54#, 8);
  gmul2_12(42) <= to_unsigned(16#56#, 8);
  gmul2_12(43) <= to_unsigned(16#58#, 8);
  gmul2_12(44) <= to_unsigned(16#5A#, 8);
  gmul2_12(45) <= to_unsigned(16#5C#, 8);
  gmul2_12(46) <= to_unsigned(16#5E#, 8);
  gmul2_12(47) <= to_unsigned(16#60#, 8);
  gmul2_12(48) <= to_unsigned(16#62#, 8);
  gmul2_12(49) <= to_unsigned(16#64#, 8);
  gmul2_12(50) <= to_unsigned(16#66#, 8);
  gmul2_12(51) <= to_unsigned(16#68#, 8);
  gmul2_12(52) <= to_unsigned(16#6A#, 8);
  gmul2_12(53) <= to_unsigned(16#6C#, 8);
  gmul2_12(54) <= to_unsigned(16#6E#, 8);
  gmul2_12(55) <= to_unsigned(16#70#, 8);
  gmul2_12(56) <= to_unsigned(16#72#, 8);
  gmul2_12(57) <= to_unsigned(16#74#, 8);
  gmul2_12(58) <= to_unsigned(16#76#, 8);
  gmul2_12(59) <= to_unsigned(16#78#, 8);
  gmul2_12(60) <= to_unsigned(16#7A#, 8);
  gmul2_12(61) <= to_unsigned(16#7C#, 8);
  gmul2_12(62) <= to_unsigned(16#7E#, 8);
  gmul2_12(63) <= to_unsigned(16#80#, 8);
  gmul2_12(64) <= to_unsigned(16#82#, 8);
  gmul2_12(65) <= to_unsigned(16#84#, 8);
  gmul2_12(66) <= to_unsigned(16#86#, 8);
  gmul2_12(67) <= to_unsigned(16#88#, 8);
  gmul2_12(68) <= to_unsigned(16#8A#, 8);
  gmul2_12(69) <= to_unsigned(16#8C#, 8);
  gmul2_12(70) <= to_unsigned(16#8E#, 8);
  gmul2_12(71) <= to_unsigned(16#90#, 8);
  gmul2_12(72) <= to_unsigned(16#92#, 8);
  gmul2_12(73) <= to_unsigned(16#94#, 8);
  gmul2_12(74) <= to_unsigned(16#96#, 8);
  gmul2_12(75) <= to_unsigned(16#98#, 8);
  gmul2_12(76) <= to_unsigned(16#9A#, 8);
  gmul2_12(77) <= to_unsigned(16#9C#, 8);
  gmul2_12(78) <= to_unsigned(16#9E#, 8);
  gmul2_12(79) <= to_unsigned(16#A0#, 8);
  gmul2_12(80) <= to_unsigned(16#A2#, 8);
  gmul2_12(81) <= to_unsigned(16#A4#, 8);
  gmul2_12(82) <= to_unsigned(16#A6#, 8);
  gmul2_12(83) <= to_unsigned(16#A8#, 8);
  gmul2_12(84) <= to_unsigned(16#AA#, 8);
  gmul2_12(85) <= to_unsigned(16#AC#, 8);
  gmul2_12(86) <= to_unsigned(16#AE#, 8);
  gmul2_12(87) <= to_unsigned(16#B0#, 8);
  gmul2_12(88) <= to_unsigned(16#B2#, 8);
  gmul2_12(89) <= to_unsigned(16#B4#, 8);
  gmul2_12(90) <= to_unsigned(16#B6#, 8);
  gmul2_12(91) <= to_unsigned(16#B8#, 8);
  gmul2_12(92) <= to_unsigned(16#BA#, 8);
  gmul2_12(93) <= to_unsigned(16#BC#, 8);
  gmul2_12(94) <= to_unsigned(16#BE#, 8);
  gmul2_12(95) <= to_unsigned(16#C0#, 8);
  gmul2_12(96) <= to_unsigned(16#C2#, 8);
  gmul2_12(97) <= to_unsigned(16#C4#, 8);
  gmul2_12(98) <= to_unsigned(16#C6#, 8);
  gmul2_12(99) <= to_unsigned(16#C8#, 8);
  gmul2_12(100) <= to_unsigned(16#CA#, 8);
  gmul2_12(101) <= to_unsigned(16#CC#, 8);
  gmul2_12(102) <= to_unsigned(16#CE#, 8);
  gmul2_12(103) <= to_unsigned(16#D0#, 8);
  gmul2_12(104) <= to_unsigned(16#D2#, 8);
  gmul2_12(105) <= to_unsigned(16#D4#, 8);
  gmul2_12(106) <= to_unsigned(16#D6#, 8);
  gmul2_12(107) <= to_unsigned(16#D8#, 8);
  gmul2_12(108) <= to_unsigned(16#DA#, 8);
  gmul2_12(109) <= to_unsigned(16#DC#, 8);
  gmul2_12(110) <= to_unsigned(16#DE#, 8);
  gmul2_12(111) <= to_unsigned(16#E0#, 8);
  gmul2_12(112) <= to_unsigned(16#E2#, 8);
  gmul2_12(113) <= to_unsigned(16#E4#, 8);
  gmul2_12(114) <= to_unsigned(16#E6#, 8);
  gmul2_12(115) <= to_unsigned(16#E8#, 8);
  gmul2_12(116) <= to_unsigned(16#EA#, 8);
  gmul2_12(117) <= to_unsigned(16#EC#, 8);
  gmul2_12(118) <= to_unsigned(16#EE#, 8);
  gmul2_12(119) <= to_unsigned(16#F0#, 8);
  gmul2_12(120) <= to_unsigned(16#F2#, 8);
  gmul2_12(121) <= to_unsigned(16#F4#, 8);
  gmul2_12(122) <= to_unsigned(16#F6#, 8);
  gmul2_12(123) <= to_unsigned(16#F8#, 8);
  gmul2_12(124) <= to_unsigned(16#FA#, 8);
  gmul2_12(125) <= to_unsigned(16#FC#, 8);
  gmul2_12(126) <= to_unsigned(16#FE#, 8);
  gmul2_12(127) <= to_unsigned(16#1B#, 8);
  gmul2_12(128) <= to_unsigned(16#19#, 8);
  gmul2_12(129) <= to_unsigned(16#1F#, 8);
  gmul2_12(130) <= to_unsigned(16#1D#, 8);
  gmul2_12(131) <= to_unsigned(16#13#, 8);
  gmul2_12(132) <= to_unsigned(16#11#, 8);
  gmul2_12(133) <= to_unsigned(16#17#, 8);
  gmul2_12(134) <= to_unsigned(16#15#, 8);
  gmul2_12(135) <= to_unsigned(16#0B#, 8);
  gmul2_12(136) <= to_unsigned(16#09#, 8);
  gmul2_12(137) <= to_unsigned(16#0F#, 8);
  gmul2_12(138) <= to_unsigned(16#0D#, 8);
  gmul2_12(139) <= to_unsigned(16#03#, 8);
  gmul2_12(140) <= to_unsigned(16#01#, 8);
  gmul2_12(141) <= to_unsigned(16#07#, 8);
  gmul2_12(142) <= to_unsigned(16#05#, 8);
  gmul2_12(143) <= to_unsigned(16#3B#, 8);
  gmul2_12(144) <= to_unsigned(16#39#, 8);
  gmul2_12(145) <= to_unsigned(16#3F#, 8);
  gmul2_12(146) <= to_unsigned(16#3D#, 8);
  gmul2_12(147) <= to_unsigned(16#33#, 8);
  gmul2_12(148) <= to_unsigned(16#31#, 8);
  gmul2_12(149) <= to_unsigned(16#37#, 8);
  gmul2_12(150) <= to_unsigned(16#35#, 8);
  gmul2_12(151) <= to_unsigned(16#2B#, 8);
  gmul2_12(152) <= to_unsigned(16#29#, 8);
  gmul2_12(153) <= to_unsigned(16#2F#, 8);
  gmul2_12(154) <= to_unsigned(16#2D#, 8);
  gmul2_12(155) <= to_unsigned(16#23#, 8);
  gmul2_12(156) <= to_unsigned(16#21#, 8);
  gmul2_12(157) <= to_unsigned(16#27#, 8);
  gmul2_12(158) <= to_unsigned(16#25#, 8);
  gmul2_12(159) <= to_unsigned(16#5B#, 8);
  gmul2_12(160) <= to_unsigned(16#59#, 8);
  gmul2_12(161) <= to_unsigned(16#5F#, 8);
  gmul2_12(162) <= to_unsigned(16#5D#, 8);
  gmul2_12(163) <= to_unsigned(16#53#, 8);
  gmul2_12(164) <= to_unsigned(16#51#, 8);
  gmul2_12(165) <= to_unsigned(16#57#, 8);
  gmul2_12(166) <= to_unsigned(16#55#, 8);
  gmul2_12(167) <= to_unsigned(16#4B#, 8);
  gmul2_12(168) <= to_unsigned(16#49#, 8);
  gmul2_12(169) <= to_unsigned(16#4F#, 8);
  gmul2_12(170) <= to_unsigned(16#4D#, 8);
  gmul2_12(171) <= to_unsigned(16#43#, 8);
  gmul2_12(172) <= to_unsigned(16#41#, 8);
  gmul2_12(173) <= to_unsigned(16#47#, 8);
  gmul2_12(174) <= to_unsigned(16#45#, 8);
  gmul2_12(175) <= to_unsigned(16#7B#, 8);
  gmul2_12(176) <= to_unsigned(16#79#, 8);
  gmul2_12(177) <= to_unsigned(16#7F#, 8);
  gmul2_12(178) <= to_unsigned(16#7D#, 8);
  gmul2_12(179) <= to_unsigned(16#73#, 8);
  gmul2_12(180) <= to_unsigned(16#71#, 8);
  gmul2_12(181) <= to_unsigned(16#77#, 8);
  gmul2_12(182) <= to_unsigned(16#75#, 8);
  gmul2_12(183) <= to_unsigned(16#6B#, 8);
  gmul2_12(184) <= to_unsigned(16#69#, 8);
  gmul2_12(185) <= to_unsigned(16#6F#, 8);
  gmul2_12(186) <= to_unsigned(16#6D#, 8);
  gmul2_12(187) <= to_unsigned(16#63#, 8);
  gmul2_12(188) <= to_unsigned(16#61#, 8);
  gmul2_12(189) <= to_unsigned(16#67#, 8);
  gmul2_12(190) <= to_unsigned(16#65#, 8);
  gmul2_12(191) <= to_unsigned(16#9B#, 8);
  gmul2_12(192) <= to_unsigned(16#99#, 8);
  gmul2_12(193) <= to_unsigned(16#9F#, 8);
  gmul2_12(194) <= to_unsigned(16#9D#, 8);
  gmul2_12(195) <= to_unsigned(16#93#, 8);
  gmul2_12(196) <= to_unsigned(16#91#, 8);
  gmul2_12(197) <= to_unsigned(16#97#, 8);
  gmul2_12(198) <= to_unsigned(16#95#, 8);
  gmul2_12(199) <= to_unsigned(16#8B#, 8);
  gmul2_12(200) <= to_unsigned(16#89#, 8);
  gmul2_12(201) <= to_unsigned(16#8F#, 8);
  gmul2_12(202) <= to_unsigned(16#8D#, 8);
  gmul2_12(203) <= to_unsigned(16#83#, 8);
  gmul2_12(204) <= to_unsigned(16#81#, 8);
  gmul2_12(205) <= to_unsigned(16#87#, 8);
  gmul2_12(206) <= to_unsigned(16#85#, 8);
  gmul2_12(207) <= to_unsigned(16#BB#, 8);
  gmul2_12(208) <= to_unsigned(16#B9#, 8);
  gmul2_12(209) <= to_unsigned(16#BF#, 8);
  gmul2_12(210) <= to_unsigned(16#BD#, 8);
  gmul2_12(211) <= to_unsigned(16#B3#, 8);
  gmul2_12(212) <= to_unsigned(16#B1#, 8);
  gmul2_12(213) <= to_unsigned(16#B7#, 8);
  gmul2_12(214) <= to_unsigned(16#B5#, 8);
  gmul2_12(215) <= to_unsigned(16#AB#, 8);
  gmul2_12(216) <= to_unsigned(16#A9#, 8);
  gmul2_12(217) <= to_unsigned(16#AF#, 8);
  gmul2_12(218) <= to_unsigned(16#AD#, 8);
  gmul2_12(219) <= to_unsigned(16#A3#, 8);
  gmul2_12(220) <= to_unsigned(16#A1#, 8);
  gmul2_12(221) <= to_unsigned(16#A7#, 8);
  gmul2_12(222) <= to_unsigned(16#A5#, 8);
  gmul2_12(223) <= to_unsigned(16#DB#, 8);
  gmul2_12(224) <= to_unsigned(16#D9#, 8);
  gmul2_12(225) <= to_unsigned(16#DF#, 8);
  gmul2_12(226) <= to_unsigned(16#DD#, 8);
  gmul2_12(227) <= to_unsigned(16#D3#, 8);
  gmul2_12(228) <= to_unsigned(16#D1#, 8);
  gmul2_12(229) <= to_unsigned(16#D7#, 8);
  gmul2_12(230) <= to_unsigned(16#D5#, 8);
  gmul2_12(231) <= to_unsigned(16#CB#, 8);
  gmul2_12(232) <= to_unsigned(16#C9#, 8);
  gmul2_12(233) <= to_unsigned(16#CF#, 8);
  gmul2_12(234) <= to_unsigned(16#CD#, 8);
  gmul2_12(235) <= to_unsigned(16#C3#, 8);
  gmul2_12(236) <= to_unsigned(16#C1#, 8);
  gmul2_12(237) <= to_unsigned(16#C7#, 8);
  gmul2_12(238) <= to_unsigned(16#C5#, 8);
  gmul2_12(239) <= to_unsigned(16#FB#, 8);
  gmul2_12(240) <= to_unsigned(16#F9#, 8);
  gmul2_12(241) <= to_unsigned(16#FF#, 8);
  gmul2_12(242) <= to_unsigned(16#FD#, 8);
  gmul2_12(243) <= to_unsigned(16#F3#, 8);
  gmul2_12(244) <= to_unsigned(16#F1#, 8);
  gmul2_12(245) <= to_unsigned(16#F7#, 8);
  gmul2_12(246) <= to_unsigned(16#F5#, 8);
  gmul2_12(247) <= to_unsigned(16#EB#, 8);
  gmul2_12(248) <= to_unsigned(16#E9#, 8);
  gmul2_12(249) <= to_unsigned(16#EF#, 8);
  gmul2_12(250) <= to_unsigned(16#ED#, 8);
  gmul2_12(251) <= to_unsigned(16#E3#, 8);
  gmul2_12(252) <= to_unsigned(16#E1#, 8);
  gmul2_12(253) <= to_unsigned(16#E7#, 8);
  gmul2_12(254) <= to_unsigned(16#E5#, 8);
  gmul2_12(255) <= to_unsigned(16#E5#, 8);

  gmul3_12(0) <= to_unsigned(16#03#, 8);
  gmul3_12(1) <= to_unsigned(16#06#, 8);
  gmul3_12(2) <= to_unsigned(16#05#, 8);
  gmul3_12(3) <= to_unsigned(16#0C#, 8);
  gmul3_12(4) <= to_unsigned(16#0F#, 8);
  gmul3_12(5) <= to_unsigned(16#0A#, 8);
  gmul3_12(6) <= to_unsigned(16#09#, 8);
  gmul3_12(7) <= to_unsigned(16#18#, 8);
  gmul3_12(8) <= to_unsigned(16#1B#, 8);
  gmul3_12(9) <= to_unsigned(16#1E#, 8);
  gmul3_12(10) <= to_unsigned(16#1D#, 8);
  gmul3_12(11) <= to_unsigned(16#14#, 8);
  gmul3_12(12) <= to_unsigned(16#17#, 8);
  gmul3_12(13) <= to_unsigned(16#12#, 8);
  gmul3_12(14) <= to_unsigned(16#11#, 8);
  gmul3_12(15) <= to_unsigned(16#30#, 8);
  gmul3_12(16) <= to_unsigned(16#33#, 8);
  gmul3_12(17) <= to_unsigned(16#36#, 8);
  gmul3_12(18) <= to_unsigned(16#35#, 8);
  gmul3_12(19) <= to_unsigned(16#3C#, 8);
  gmul3_12(20) <= to_unsigned(16#3F#, 8);
  gmul3_12(21) <= to_unsigned(16#3A#, 8);
  gmul3_12(22) <= to_unsigned(16#39#, 8);
  gmul3_12(23) <= to_unsigned(16#28#, 8);
  gmul3_12(24) <= to_unsigned(16#2B#, 8);
  gmul3_12(25) <= to_unsigned(16#2E#, 8);
  gmul3_12(26) <= to_unsigned(16#2D#, 8);
  gmul3_12(27) <= to_unsigned(16#24#, 8);
  gmul3_12(28) <= to_unsigned(16#27#, 8);
  gmul3_12(29) <= to_unsigned(16#22#, 8);
  gmul3_12(30) <= to_unsigned(16#21#, 8);
  gmul3_12(31) <= to_unsigned(16#60#, 8);
  gmul3_12(32) <= to_unsigned(16#63#, 8);
  gmul3_12(33) <= to_unsigned(16#66#, 8);
  gmul3_12(34) <= to_unsigned(16#65#, 8);
  gmul3_12(35) <= to_unsigned(16#6C#, 8);
  gmul3_12(36) <= to_unsigned(16#6F#, 8);
  gmul3_12(37) <= to_unsigned(16#6A#, 8);
  gmul3_12(38) <= to_unsigned(16#69#, 8);
  gmul3_12(39) <= to_unsigned(16#78#, 8);
  gmul3_12(40) <= to_unsigned(16#7B#, 8);
  gmul3_12(41) <= to_unsigned(16#7E#, 8);
  gmul3_12(42) <= to_unsigned(16#7D#, 8);
  gmul3_12(43) <= to_unsigned(16#74#, 8);
  gmul3_12(44) <= to_unsigned(16#77#, 8);
  gmul3_12(45) <= to_unsigned(16#72#, 8);
  gmul3_12(46) <= to_unsigned(16#71#, 8);
  gmul3_12(47) <= to_unsigned(16#50#, 8);
  gmul3_12(48) <= to_unsigned(16#53#, 8);
  gmul3_12(49) <= to_unsigned(16#56#, 8);
  gmul3_12(50) <= to_unsigned(16#55#, 8);
  gmul3_12(51) <= to_unsigned(16#5C#, 8);
  gmul3_12(52) <= to_unsigned(16#5F#, 8);
  gmul3_12(53) <= to_unsigned(16#5A#, 8);
  gmul3_12(54) <= to_unsigned(16#59#, 8);
  gmul3_12(55) <= to_unsigned(16#48#, 8);
  gmul3_12(56) <= to_unsigned(16#4B#, 8);
  gmul3_12(57) <= to_unsigned(16#4E#, 8);
  gmul3_12(58) <= to_unsigned(16#4D#, 8);
  gmul3_12(59) <= to_unsigned(16#44#, 8);
  gmul3_12(60) <= to_unsigned(16#47#, 8);
  gmul3_12(61) <= to_unsigned(16#42#, 8);
  gmul3_12(62) <= to_unsigned(16#41#, 8);
  gmul3_12(63) <= to_unsigned(16#C0#, 8);
  gmul3_12(64) <= to_unsigned(16#C3#, 8);
  gmul3_12(65) <= to_unsigned(16#C6#, 8);
  gmul3_12(66) <= to_unsigned(16#C5#, 8);
  gmul3_12(67) <= to_unsigned(16#CC#, 8);
  gmul3_12(68) <= to_unsigned(16#CF#, 8);
  gmul3_12(69) <= to_unsigned(16#CA#, 8);
  gmul3_12(70) <= to_unsigned(16#C9#, 8);
  gmul3_12(71) <= to_unsigned(16#D8#, 8);
  gmul3_12(72) <= to_unsigned(16#DB#, 8);
  gmul3_12(73) <= to_unsigned(16#DE#, 8);
  gmul3_12(74) <= to_unsigned(16#DD#, 8);
  gmul3_12(75) <= to_unsigned(16#D4#, 8);
  gmul3_12(76) <= to_unsigned(16#D7#, 8);
  gmul3_12(77) <= to_unsigned(16#D2#, 8);
  gmul3_12(78) <= to_unsigned(16#D1#, 8);
  gmul3_12(79) <= to_unsigned(16#F0#, 8);
  gmul3_12(80) <= to_unsigned(16#F3#, 8);
  gmul3_12(81) <= to_unsigned(16#F6#, 8);
  gmul3_12(82) <= to_unsigned(16#F5#, 8);
  gmul3_12(83) <= to_unsigned(16#FC#, 8);
  gmul3_12(84) <= to_unsigned(16#FF#, 8);
  gmul3_12(85) <= to_unsigned(16#FA#, 8);
  gmul3_12(86) <= to_unsigned(16#F9#, 8);
  gmul3_12(87) <= to_unsigned(16#E8#, 8);
  gmul3_12(88) <= to_unsigned(16#EB#, 8);
  gmul3_12(89) <= to_unsigned(16#EE#, 8);
  gmul3_12(90) <= to_unsigned(16#ED#, 8);
  gmul3_12(91) <= to_unsigned(16#E4#, 8);
  gmul3_12(92) <= to_unsigned(16#E7#, 8);
  gmul3_12(93) <= to_unsigned(16#E2#, 8);
  gmul3_12(94) <= to_unsigned(16#E1#, 8);
  gmul3_12(95) <= to_unsigned(16#A0#, 8);
  gmul3_12(96) <= to_unsigned(16#A3#, 8);
  gmul3_12(97) <= to_unsigned(16#A6#, 8);
  gmul3_12(98) <= to_unsigned(16#A5#, 8);
  gmul3_12(99) <= to_unsigned(16#AC#, 8);
  gmul3_12(100) <= to_unsigned(16#AF#, 8);
  gmul3_12(101) <= to_unsigned(16#AA#, 8);
  gmul3_12(102) <= to_unsigned(16#A9#, 8);
  gmul3_12(103) <= to_unsigned(16#B8#, 8);
  gmul3_12(104) <= to_unsigned(16#BB#, 8);
  gmul3_12(105) <= to_unsigned(16#BE#, 8);
  gmul3_12(106) <= to_unsigned(16#BD#, 8);
  gmul3_12(107) <= to_unsigned(16#B4#, 8);
  gmul3_12(108) <= to_unsigned(16#B7#, 8);
  gmul3_12(109) <= to_unsigned(16#B2#, 8);
  gmul3_12(110) <= to_unsigned(16#B1#, 8);
  gmul3_12(111) <= to_unsigned(16#90#, 8);
  gmul3_12(112) <= to_unsigned(16#93#, 8);
  gmul3_12(113) <= to_unsigned(16#96#, 8);
  gmul3_12(114) <= to_unsigned(16#95#, 8);
  gmul3_12(115) <= to_unsigned(16#9C#, 8);
  gmul3_12(116) <= to_unsigned(16#9F#, 8);
  gmul3_12(117) <= to_unsigned(16#9A#, 8);
  gmul3_12(118) <= to_unsigned(16#99#, 8);
  gmul3_12(119) <= to_unsigned(16#88#, 8);
  gmul3_12(120) <= to_unsigned(16#8B#, 8);
  gmul3_12(121) <= to_unsigned(16#8E#, 8);
  gmul3_12(122) <= to_unsigned(16#8D#, 8);
  gmul3_12(123) <= to_unsigned(16#84#, 8);
  gmul3_12(124) <= to_unsigned(16#87#, 8);
  gmul3_12(125) <= to_unsigned(16#82#, 8);
  gmul3_12(126) <= to_unsigned(16#81#, 8);
  gmul3_12(127) <= to_unsigned(16#9B#, 8);
  gmul3_12(128) <= to_unsigned(16#98#, 8);
  gmul3_12(129) <= to_unsigned(16#9D#, 8);
  gmul3_12(130) <= to_unsigned(16#9E#, 8);
  gmul3_12(131) <= to_unsigned(16#97#, 8);
  gmul3_12(132) <= to_unsigned(16#94#, 8);
  gmul3_12(133) <= to_unsigned(16#91#, 8);
  gmul3_12(134) <= to_unsigned(16#92#, 8);
  gmul3_12(135) <= to_unsigned(16#83#, 8);
  gmul3_12(136) <= to_unsigned(16#80#, 8);
  gmul3_12(137) <= to_unsigned(16#85#, 8);
  gmul3_12(138) <= to_unsigned(16#86#, 8);
  gmul3_12(139) <= to_unsigned(16#8F#, 8);
  gmul3_12(140) <= to_unsigned(16#8C#, 8);
  gmul3_12(141) <= to_unsigned(16#89#, 8);
  gmul3_12(142) <= to_unsigned(16#8A#, 8);
  gmul3_12(143) <= to_unsigned(16#AB#, 8);
  gmul3_12(144) <= to_unsigned(16#A8#, 8);
  gmul3_12(145) <= to_unsigned(16#AD#, 8);
  gmul3_12(146) <= to_unsigned(16#AE#, 8);
  gmul3_12(147) <= to_unsigned(16#A7#, 8);
  gmul3_12(148) <= to_unsigned(16#A4#, 8);
  gmul3_12(149) <= to_unsigned(16#A1#, 8);
  gmul3_12(150) <= to_unsigned(16#A2#, 8);
  gmul3_12(151) <= to_unsigned(16#B3#, 8);
  gmul3_12(152) <= to_unsigned(16#B0#, 8);
  gmul3_12(153) <= to_unsigned(16#B5#, 8);
  gmul3_12(154) <= to_unsigned(16#B6#, 8);
  gmul3_12(155) <= to_unsigned(16#BF#, 8);
  gmul3_12(156) <= to_unsigned(16#BC#, 8);
  gmul3_12(157) <= to_unsigned(16#B9#, 8);
  gmul3_12(158) <= to_unsigned(16#BA#, 8);
  gmul3_12(159) <= to_unsigned(16#FB#, 8);
  gmul3_12(160) <= to_unsigned(16#F8#, 8);
  gmul3_12(161) <= to_unsigned(16#FD#, 8);
  gmul3_12(162) <= to_unsigned(16#FE#, 8);
  gmul3_12(163) <= to_unsigned(16#F7#, 8);
  gmul3_12(164) <= to_unsigned(16#F4#, 8);
  gmul3_12(165) <= to_unsigned(16#F1#, 8);
  gmul3_12(166) <= to_unsigned(16#F2#, 8);
  gmul3_12(167) <= to_unsigned(16#E3#, 8);
  gmul3_12(168) <= to_unsigned(16#E0#, 8);
  gmul3_12(169) <= to_unsigned(16#E5#, 8);
  gmul3_12(170) <= to_unsigned(16#E6#, 8);
  gmul3_12(171) <= to_unsigned(16#EF#, 8);
  gmul3_12(172) <= to_unsigned(16#EC#, 8);
  gmul3_12(173) <= to_unsigned(16#E9#, 8);
  gmul3_12(174) <= to_unsigned(16#EA#, 8);
  gmul3_12(175) <= to_unsigned(16#CB#, 8);
  gmul3_12(176) <= to_unsigned(16#C8#, 8);
  gmul3_12(177) <= to_unsigned(16#CD#, 8);
  gmul3_12(178) <= to_unsigned(16#CE#, 8);
  gmul3_12(179) <= to_unsigned(16#C7#, 8);
  gmul3_12(180) <= to_unsigned(16#C4#, 8);
  gmul3_12(181) <= to_unsigned(16#C1#, 8);
  gmul3_12(182) <= to_unsigned(16#C2#, 8);
  gmul3_12(183) <= to_unsigned(16#D3#, 8);
  gmul3_12(184) <= to_unsigned(16#D0#, 8);
  gmul3_12(185) <= to_unsigned(16#D5#, 8);
  gmul3_12(186) <= to_unsigned(16#D6#, 8);
  gmul3_12(187) <= to_unsigned(16#DF#, 8);
  gmul3_12(188) <= to_unsigned(16#DC#, 8);
  gmul3_12(189) <= to_unsigned(16#D9#, 8);
  gmul3_12(190) <= to_unsigned(16#DA#, 8);
  gmul3_12(191) <= to_unsigned(16#5B#, 8);
  gmul3_12(192) <= to_unsigned(16#58#, 8);
  gmul3_12(193) <= to_unsigned(16#5D#, 8);
  gmul3_12(194) <= to_unsigned(16#5E#, 8);
  gmul3_12(195) <= to_unsigned(16#57#, 8);
  gmul3_12(196) <= to_unsigned(16#54#, 8);
  gmul3_12(197) <= to_unsigned(16#51#, 8);
  gmul3_12(198) <= to_unsigned(16#52#, 8);
  gmul3_12(199) <= to_unsigned(16#43#, 8);
  gmul3_12(200) <= to_unsigned(16#40#, 8);
  gmul3_12(201) <= to_unsigned(16#45#, 8);
  gmul3_12(202) <= to_unsigned(16#46#, 8);
  gmul3_12(203) <= to_unsigned(16#4F#, 8);
  gmul3_12(204) <= to_unsigned(16#4C#, 8);
  gmul3_12(205) <= to_unsigned(16#49#, 8);
  gmul3_12(206) <= to_unsigned(16#4A#, 8);
  gmul3_12(207) <= to_unsigned(16#6B#, 8);
  gmul3_12(208) <= to_unsigned(16#68#, 8);
  gmul3_12(209) <= to_unsigned(16#6D#, 8);
  gmul3_12(210) <= to_unsigned(16#6E#, 8);
  gmul3_12(211) <= to_unsigned(16#67#, 8);
  gmul3_12(212) <= to_unsigned(16#64#, 8);
  gmul3_12(213) <= to_unsigned(16#61#, 8);
  gmul3_12(214) <= to_unsigned(16#62#, 8);
  gmul3_12(215) <= to_unsigned(16#73#, 8);
  gmul3_12(216) <= to_unsigned(16#70#, 8);
  gmul3_12(217) <= to_unsigned(16#75#, 8);
  gmul3_12(218) <= to_unsigned(16#76#, 8);
  gmul3_12(219) <= to_unsigned(16#7F#, 8);
  gmul3_12(220) <= to_unsigned(16#7C#, 8);
  gmul3_12(221) <= to_unsigned(16#79#, 8);
  gmul3_12(222) <= to_unsigned(16#7A#, 8);
  gmul3_12(223) <= to_unsigned(16#3B#, 8);
  gmul3_12(224) <= to_unsigned(16#38#, 8);
  gmul3_12(225) <= to_unsigned(16#3D#, 8);
  gmul3_12(226) <= to_unsigned(16#3E#, 8);
  gmul3_12(227) <= to_unsigned(16#37#, 8);
  gmul3_12(228) <= to_unsigned(16#34#, 8);
  gmul3_12(229) <= to_unsigned(16#31#, 8);
  gmul3_12(230) <= to_unsigned(16#32#, 8);
  gmul3_12(231) <= to_unsigned(16#23#, 8);
  gmul3_12(232) <= to_unsigned(16#20#, 8);
  gmul3_12(233) <= to_unsigned(16#25#, 8);
  gmul3_12(234) <= to_unsigned(16#26#, 8);
  gmul3_12(235) <= to_unsigned(16#2F#, 8);
  gmul3_12(236) <= to_unsigned(16#2C#, 8);
  gmul3_12(237) <= to_unsigned(16#29#, 8);
  gmul3_12(238) <= to_unsigned(16#2A#, 8);
  gmul3_12(239) <= to_unsigned(16#0B#, 8);
  gmul3_12(240) <= to_unsigned(16#08#, 8);
  gmul3_12(241) <= to_unsigned(16#0D#, 8);
  gmul3_12(242) <= to_unsigned(16#0E#, 8);
  gmul3_12(243) <= to_unsigned(16#07#, 8);
  gmul3_12(244) <= to_unsigned(16#04#, 8);
  gmul3_12(245) <= to_unsigned(16#01#, 8);
  gmul3_12(246) <= to_unsigned(16#02#, 8);
  gmul3_12(247) <= to_unsigned(16#13#, 8);
  gmul3_12(248) <= to_unsigned(16#10#, 8);
  gmul3_12(249) <= to_unsigned(16#15#, 8);
  gmul3_12(250) <= to_unsigned(16#16#, 8);
  gmul3_12(251) <= to_unsigned(16#1F#, 8);
  gmul3_12(252) <= to_unsigned(16#1C#, 8);
  gmul3_12(253) <= to_unsigned(16#19#, 8);
  gmul3_12(254) <= to_unsigned(16#1A#, 8);
  gmul3_12(255) <= to_unsigned(16#1A#, 8);

  gmul2_13(0) <= to_unsigned(16#02#, 8);
  gmul2_13(1) <= to_unsigned(16#04#, 8);
  gmul2_13(2) <= to_unsigned(16#06#, 8);
  gmul2_13(3) <= to_unsigned(16#08#, 8);
  gmul2_13(4) <= to_unsigned(16#0A#, 8);
  gmul2_13(5) <= to_unsigned(16#0C#, 8);
  gmul2_13(6) <= to_unsigned(16#0E#, 8);
  gmul2_13(7) <= to_unsigned(16#10#, 8);
  gmul2_13(8) <= to_unsigned(16#12#, 8);
  gmul2_13(9) <= to_unsigned(16#14#, 8);
  gmul2_13(10) <= to_unsigned(16#16#, 8);
  gmul2_13(11) <= to_unsigned(16#18#, 8);
  gmul2_13(12) <= to_unsigned(16#1A#, 8);
  gmul2_13(13) <= to_unsigned(16#1C#, 8);
  gmul2_13(14) <= to_unsigned(16#1E#, 8);
  gmul2_13(15) <= to_unsigned(16#20#, 8);
  gmul2_13(16) <= to_unsigned(16#22#, 8);
  gmul2_13(17) <= to_unsigned(16#24#, 8);
  gmul2_13(18) <= to_unsigned(16#26#, 8);
  gmul2_13(19) <= to_unsigned(16#28#, 8);
  gmul2_13(20) <= to_unsigned(16#2A#, 8);
  gmul2_13(21) <= to_unsigned(16#2C#, 8);
  gmul2_13(22) <= to_unsigned(16#2E#, 8);
  gmul2_13(23) <= to_unsigned(16#30#, 8);
  gmul2_13(24) <= to_unsigned(16#32#, 8);
  gmul2_13(25) <= to_unsigned(16#34#, 8);
  gmul2_13(26) <= to_unsigned(16#36#, 8);
  gmul2_13(27) <= to_unsigned(16#38#, 8);
  gmul2_13(28) <= to_unsigned(16#3A#, 8);
  gmul2_13(29) <= to_unsigned(16#3C#, 8);
  gmul2_13(30) <= to_unsigned(16#3E#, 8);
  gmul2_13(31) <= to_unsigned(16#40#, 8);
  gmul2_13(32) <= to_unsigned(16#42#, 8);
  gmul2_13(33) <= to_unsigned(16#44#, 8);
  gmul2_13(34) <= to_unsigned(16#46#, 8);
  gmul2_13(35) <= to_unsigned(16#48#, 8);
  gmul2_13(36) <= to_unsigned(16#4A#, 8);
  gmul2_13(37) <= to_unsigned(16#4C#, 8);
  gmul2_13(38) <= to_unsigned(16#4E#, 8);
  gmul2_13(39) <= to_unsigned(16#50#, 8);
  gmul2_13(40) <= to_unsigned(16#52#, 8);
  gmul2_13(41) <= to_unsigned(16#54#, 8);
  gmul2_13(42) <= to_unsigned(16#56#, 8);
  gmul2_13(43) <= to_unsigned(16#58#, 8);
  gmul2_13(44) <= to_unsigned(16#5A#, 8);
  gmul2_13(45) <= to_unsigned(16#5C#, 8);
  gmul2_13(46) <= to_unsigned(16#5E#, 8);
  gmul2_13(47) <= to_unsigned(16#60#, 8);
  gmul2_13(48) <= to_unsigned(16#62#, 8);
  gmul2_13(49) <= to_unsigned(16#64#, 8);
  gmul2_13(50) <= to_unsigned(16#66#, 8);
  gmul2_13(51) <= to_unsigned(16#68#, 8);
  gmul2_13(52) <= to_unsigned(16#6A#, 8);
  gmul2_13(53) <= to_unsigned(16#6C#, 8);
  gmul2_13(54) <= to_unsigned(16#6E#, 8);
  gmul2_13(55) <= to_unsigned(16#70#, 8);
  gmul2_13(56) <= to_unsigned(16#72#, 8);
  gmul2_13(57) <= to_unsigned(16#74#, 8);
  gmul2_13(58) <= to_unsigned(16#76#, 8);
  gmul2_13(59) <= to_unsigned(16#78#, 8);
  gmul2_13(60) <= to_unsigned(16#7A#, 8);
  gmul2_13(61) <= to_unsigned(16#7C#, 8);
  gmul2_13(62) <= to_unsigned(16#7E#, 8);
  gmul2_13(63) <= to_unsigned(16#80#, 8);
  gmul2_13(64) <= to_unsigned(16#82#, 8);
  gmul2_13(65) <= to_unsigned(16#84#, 8);
  gmul2_13(66) <= to_unsigned(16#86#, 8);
  gmul2_13(67) <= to_unsigned(16#88#, 8);
  gmul2_13(68) <= to_unsigned(16#8A#, 8);
  gmul2_13(69) <= to_unsigned(16#8C#, 8);
  gmul2_13(70) <= to_unsigned(16#8E#, 8);
  gmul2_13(71) <= to_unsigned(16#90#, 8);
  gmul2_13(72) <= to_unsigned(16#92#, 8);
  gmul2_13(73) <= to_unsigned(16#94#, 8);
  gmul2_13(74) <= to_unsigned(16#96#, 8);
  gmul2_13(75) <= to_unsigned(16#98#, 8);
  gmul2_13(76) <= to_unsigned(16#9A#, 8);
  gmul2_13(77) <= to_unsigned(16#9C#, 8);
  gmul2_13(78) <= to_unsigned(16#9E#, 8);
  gmul2_13(79) <= to_unsigned(16#A0#, 8);
  gmul2_13(80) <= to_unsigned(16#A2#, 8);
  gmul2_13(81) <= to_unsigned(16#A4#, 8);
  gmul2_13(82) <= to_unsigned(16#A6#, 8);
  gmul2_13(83) <= to_unsigned(16#A8#, 8);
  gmul2_13(84) <= to_unsigned(16#AA#, 8);
  gmul2_13(85) <= to_unsigned(16#AC#, 8);
  gmul2_13(86) <= to_unsigned(16#AE#, 8);
  gmul2_13(87) <= to_unsigned(16#B0#, 8);
  gmul2_13(88) <= to_unsigned(16#B2#, 8);
  gmul2_13(89) <= to_unsigned(16#B4#, 8);
  gmul2_13(90) <= to_unsigned(16#B6#, 8);
  gmul2_13(91) <= to_unsigned(16#B8#, 8);
  gmul2_13(92) <= to_unsigned(16#BA#, 8);
  gmul2_13(93) <= to_unsigned(16#BC#, 8);
  gmul2_13(94) <= to_unsigned(16#BE#, 8);
  gmul2_13(95) <= to_unsigned(16#C0#, 8);
  gmul2_13(96) <= to_unsigned(16#C2#, 8);
  gmul2_13(97) <= to_unsigned(16#C4#, 8);
  gmul2_13(98) <= to_unsigned(16#C6#, 8);
  gmul2_13(99) <= to_unsigned(16#C8#, 8);
  gmul2_13(100) <= to_unsigned(16#CA#, 8);
  gmul2_13(101) <= to_unsigned(16#CC#, 8);
  gmul2_13(102) <= to_unsigned(16#CE#, 8);
  gmul2_13(103) <= to_unsigned(16#D0#, 8);
  gmul2_13(104) <= to_unsigned(16#D2#, 8);
  gmul2_13(105) <= to_unsigned(16#D4#, 8);
  gmul2_13(106) <= to_unsigned(16#D6#, 8);
  gmul2_13(107) <= to_unsigned(16#D8#, 8);
  gmul2_13(108) <= to_unsigned(16#DA#, 8);
  gmul2_13(109) <= to_unsigned(16#DC#, 8);
  gmul2_13(110) <= to_unsigned(16#DE#, 8);
  gmul2_13(111) <= to_unsigned(16#E0#, 8);
  gmul2_13(112) <= to_unsigned(16#E2#, 8);
  gmul2_13(113) <= to_unsigned(16#E4#, 8);
  gmul2_13(114) <= to_unsigned(16#E6#, 8);
  gmul2_13(115) <= to_unsigned(16#E8#, 8);
  gmul2_13(116) <= to_unsigned(16#EA#, 8);
  gmul2_13(117) <= to_unsigned(16#EC#, 8);
  gmul2_13(118) <= to_unsigned(16#EE#, 8);
  gmul2_13(119) <= to_unsigned(16#F0#, 8);
  gmul2_13(120) <= to_unsigned(16#F2#, 8);
  gmul2_13(121) <= to_unsigned(16#F4#, 8);
  gmul2_13(122) <= to_unsigned(16#F6#, 8);
  gmul2_13(123) <= to_unsigned(16#F8#, 8);
  gmul2_13(124) <= to_unsigned(16#FA#, 8);
  gmul2_13(125) <= to_unsigned(16#FC#, 8);
  gmul2_13(126) <= to_unsigned(16#FE#, 8);
  gmul2_13(127) <= to_unsigned(16#1B#, 8);
  gmul2_13(128) <= to_unsigned(16#19#, 8);
  gmul2_13(129) <= to_unsigned(16#1F#, 8);
  gmul2_13(130) <= to_unsigned(16#1D#, 8);
  gmul2_13(131) <= to_unsigned(16#13#, 8);
  gmul2_13(132) <= to_unsigned(16#11#, 8);
  gmul2_13(133) <= to_unsigned(16#17#, 8);
  gmul2_13(134) <= to_unsigned(16#15#, 8);
  gmul2_13(135) <= to_unsigned(16#0B#, 8);
  gmul2_13(136) <= to_unsigned(16#09#, 8);
  gmul2_13(137) <= to_unsigned(16#0F#, 8);
  gmul2_13(138) <= to_unsigned(16#0D#, 8);
  gmul2_13(139) <= to_unsigned(16#03#, 8);
  gmul2_13(140) <= to_unsigned(16#01#, 8);
  gmul2_13(141) <= to_unsigned(16#07#, 8);
  gmul2_13(142) <= to_unsigned(16#05#, 8);
  gmul2_13(143) <= to_unsigned(16#3B#, 8);
  gmul2_13(144) <= to_unsigned(16#39#, 8);
  gmul2_13(145) <= to_unsigned(16#3F#, 8);
  gmul2_13(146) <= to_unsigned(16#3D#, 8);
  gmul2_13(147) <= to_unsigned(16#33#, 8);
  gmul2_13(148) <= to_unsigned(16#31#, 8);
  gmul2_13(149) <= to_unsigned(16#37#, 8);
  gmul2_13(150) <= to_unsigned(16#35#, 8);
  gmul2_13(151) <= to_unsigned(16#2B#, 8);
  gmul2_13(152) <= to_unsigned(16#29#, 8);
  gmul2_13(153) <= to_unsigned(16#2F#, 8);
  gmul2_13(154) <= to_unsigned(16#2D#, 8);
  gmul2_13(155) <= to_unsigned(16#23#, 8);
  gmul2_13(156) <= to_unsigned(16#21#, 8);
  gmul2_13(157) <= to_unsigned(16#27#, 8);
  gmul2_13(158) <= to_unsigned(16#25#, 8);
  gmul2_13(159) <= to_unsigned(16#5B#, 8);
  gmul2_13(160) <= to_unsigned(16#59#, 8);
  gmul2_13(161) <= to_unsigned(16#5F#, 8);
  gmul2_13(162) <= to_unsigned(16#5D#, 8);
  gmul2_13(163) <= to_unsigned(16#53#, 8);
  gmul2_13(164) <= to_unsigned(16#51#, 8);
  gmul2_13(165) <= to_unsigned(16#57#, 8);
  gmul2_13(166) <= to_unsigned(16#55#, 8);
  gmul2_13(167) <= to_unsigned(16#4B#, 8);
  gmul2_13(168) <= to_unsigned(16#49#, 8);
  gmul2_13(169) <= to_unsigned(16#4F#, 8);
  gmul2_13(170) <= to_unsigned(16#4D#, 8);
  gmul2_13(171) <= to_unsigned(16#43#, 8);
  gmul2_13(172) <= to_unsigned(16#41#, 8);
  gmul2_13(173) <= to_unsigned(16#47#, 8);
  gmul2_13(174) <= to_unsigned(16#45#, 8);
  gmul2_13(175) <= to_unsigned(16#7B#, 8);
  gmul2_13(176) <= to_unsigned(16#79#, 8);
  gmul2_13(177) <= to_unsigned(16#7F#, 8);
  gmul2_13(178) <= to_unsigned(16#7D#, 8);
  gmul2_13(179) <= to_unsigned(16#73#, 8);
  gmul2_13(180) <= to_unsigned(16#71#, 8);
  gmul2_13(181) <= to_unsigned(16#77#, 8);
  gmul2_13(182) <= to_unsigned(16#75#, 8);
  gmul2_13(183) <= to_unsigned(16#6B#, 8);
  gmul2_13(184) <= to_unsigned(16#69#, 8);
  gmul2_13(185) <= to_unsigned(16#6F#, 8);
  gmul2_13(186) <= to_unsigned(16#6D#, 8);
  gmul2_13(187) <= to_unsigned(16#63#, 8);
  gmul2_13(188) <= to_unsigned(16#61#, 8);
  gmul2_13(189) <= to_unsigned(16#67#, 8);
  gmul2_13(190) <= to_unsigned(16#65#, 8);
  gmul2_13(191) <= to_unsigned(16#9B#, 8);
  gmul2_13(192) <= to_unsigned(16#99#, 8);
  gmul2_13(193) <= to_unsigned(16#9F#, 8);
  gmul2_13(194) <= to_unsigned(16#9D#, 8);
  gmul2_13(195) <= to_unsigned(16#93#, 8);
  gmul2_13(196) <= to_unsigned(16#91#, 8);
  gmul2_13(197) <= to_unsigned(16#97#, 8);
  gmul2_13(198) <= to_unsigned(16#95#, 8);
  gmul2_13(199) <= to_unsigned(16#8B#, 8);
  gmul2_13(200) <= to_unsigned(16#89#, 8);
  gmul2_13(201) <= to_unsigned(16#8F#, 8);
  gmul2_13(202) <= to_unsigned(16#8D#, 8);
  gmul2_13(203) <= to_unsigned(16#83#, 8);
  gmul2_13(204) <= to_unsigned(16#81#, 8);
  gmul2_13(205) <= to_unsigned(16#87#, 8);
  gmul2_13(206) <= to_unsigned(16#85#, 8);
  gmul2_13(207) <= to_unsigned(16#BB#, 8);
  gmul2_13(208) <= to_unsigned(16#B9#, 8);
  gmul2_13(209) <= to_unsigned(16#BF#, 8);
  gmul2_13(210) <= to_unsigned(16#BD#, 8);
  gmul2_13(211) <= to_unsigned(16#B3#, 8);
  gmul2_13(212) <= to_unsigned(16#B1#, 8);
  gmul2_13(213) <= to_unsigned(16#B7#, 8);
  gmul2_13(214) <= to_unsigned(16#B5#, 8);
  gmul2_13(215) <= to_unsigned(16#AB#, 8);
  gmul2_13(216) <= to_unsigned(16#A9#, 8);
  gmul2_13(217) <= to_unsigned(16#AF#, 8);
  gmul2_13(218) <= to_unsigned(16#AD#, 8);
  gmul2_13(219) <= to_unsigned(16#A3#, 8);
  gmul2_13(220) <= to_unsigned(16#A1#, 8);
  gmul2_13(221) <= to_unsigned(16#A7#, 8);
  gmul2_13(222) <= to_unsigned(16#A5#, 8);
  gmul2_13(223) <= to_unsigned(16#DB#, 8);
  gmul2_13(224) <= to_unsigned(16#D9#, 8);
  gmul2_13(225) <= to_unsigned(16#DF#, 8);
  gmul2_13(226) <= to_unsigned(16#DD#, 8);
  gmul2_13(227) <= to_unsigned(16#D3#, 8);
  gmul2_13(228) <= to_unsigned(16#D1#, 8);
  gmul2_13(229) <= to_unsigned(16#D7#, 8);
  gmul2_13(230) <= to_unsigned(16#D5#, 8);
  gmul2_13(231) <= to_unsigned(16#CB#, 8);
  gmul2_13(232) <= to_unsigned(16#C9#, 8);
  gmul2_13(233) <= to_unsigned(16#CF#, 8);
  gmul2_13(234) <= to_unsigned(16#CD#, 8);
  gmul2_13(235) <= to_unsigned(16#C3#, 8);
  gmul2_13(236) <= to_unsigned(16#C1#, 8);
  gmul2_13(237) <= to_unsigned(16#C7#, 8);
  gmul2_13(238) <= to_unsigned(16#C5#, 8);
  gmul2_13(239) <= to_unsigned(16#FB#, 8);
  gmul2_13(240) <= to_unsigned(16#F9#, 8);
  gmul2_13(241) <= to_unsigned(16#FF#, 8);
  gmul2_13(242) <= to_unsigned(16#FD#, 8);
  gmul2_13(243) <= to_unsigned(16#F3#, 8);
  gmul2_13(244) <= to_unsigned(16#F1#, 8);
  gmul2_13(245) <= to_unsigned(16#F7#, 8);
  gmul2_13(246) <= to_unsigned(16#F5#, 8);
  gmul2_13(247) <= to_unsigned(16#EB#, 8);
  gmul2_13(248) <= to_unsigned(16#E9#, 8);
  gmul2_13(249) <= to_unsigned(16#EF#, 8);
  gmul2_13(250) <= to_unsigned(16#ED#, 8);
  gmul2_13(251) <= to_unsigned(16#E3#, 8);
  gmul2_13(252) <= to_unsigned(16#E1#, 8);
  gmul2_13(253) <= to_unsigned(16#E7#, 8);
  gmul2_13(254) <= to_unsigned(16#E5#, 8);
  gmul2_13(255) <= to_unsigned(16#E5#, 8);

  gmul3_13(0) <= to_unsigned(16#03#, 8);
  gmul3_13(1) <= to_unsigned(16#06#, 8);
  gmul3_13(2) <= to_unsigned(16#05#, 8);
  gmul3_13(3) <= to_unsigned(16#0C#, 8);
  gmul3_13(4) <= to_unsigned(16#0F#, 8);
  gmul3_13(5) <= to_unsigned(16#0A#, 8);
  gmul3_13(6) <= to_unsigned(16#09#, 8);
  gmul3_13(7) <= to_unsigned(16#18#, 8);
  gmul3_13(8) <= to_unsigned(16#1B#, 8);
  gmul3_13(9) <= to_unsigned(16#1E#, 8);
  gmul3_13(10) <= to_unsigned(16#1D#, 8);
  gmul3_13(11) <= to_unsigned(16#14#, 8);
  gmul3_13(12) <= to_unsigned(16#17#, 8);
  gmul3_13(13) <= to_unsigned(16#12#, 8);
  gmul3_13(14) <= to_unsigned(16#11#, 8);
  gmul3_13(15) <= to_unsigned(16#30#, 8);
  gmul3_13(16) <= to_unsigned(16#33#, 8);
  gmul3_13(17) <= to_unsigned(16#36#, 8);
  gmul3_13(18) <= to_unsigned(16#35#, 8);
  gmul3_13(19) <= to_unsigned(16#3C#, 8);
  gmul3_13(20) <= to_unsigned(16#3F#, 8);
  gmul3_13(21) <= to_unsigned(16#3A#, 8);
  gmul3_13(22) <= to_unsigned(16#39#, 8);
  gmul3_13(23) <= to_unsigned(16#28#, 8);
  gmul3_13(24) <= to_unsigned(16#2B#, 8);
  gmul3_13(25) <= to_unsigned(16#2E#, 8);
  gmul3_13(26) <= to_unsigned(16#2D#, 8);
  gmul3_13(27) <= to_unsigned(16#24#, 8);
  gmul3_13(28) <= to_unsigned(16#27#, 8);
  gmul3_13(29) <= to_unsigned(16#22#, 8);
  gmul3_13(30) <= to_unsigned(16#21#, 8);
  gmul3_13(31) <= to_unsigned(16#60#, 8);
  gmul3_13(32) <= to_unsigned(16#63#, 8);
  gmul3_13(33) <= to_unsigned(16#66#, 8);
  gmul3_13(34) <= to_unsigned(16#65#, 8);
  gmul3_13(35) <= to_unsigned(16#6C#, 8);
  gmul3_13(36) <= to_unsigned(16#6F#, 8);
  gmul3_13(37) <= to_unsigned(16#6A#, 8);
  gmul3_13(38) <= to_unsigned(16#69#, 8);
  gmul3_13(39) <= to_unsigned(16#78#, 8);
  gmul3_13(40) <= to_unsigned(16#7B#, 8);
  gmul3_13(41) <= to_unsigned(16#7E#, 8);
  gmul3_13(42) <= to_unsigned(16#7D#, 8);
  gmul3_13(43) <= to_unsigned(16#74#, 8);
  gmul3_13(44) <= to_unsigned(16#77#, 8);
  gmul3_13(45) <= to_unsigned(16#72#, 8);
  gmul3_13(46) <= to_unsigned(16#71#, 8);
  gmul3_13(47) <= to_unsigned(16#50#, 8);
  gmul3_13(48) <= to_unsigned(16#53#, 8);
  gmul3_13(49) <= to_unsigned(16#56#, 8);
  gmul3_13(50) <= to_unsigned(16#55#, 8);
  gmul3_13(51) <= to_unsigned(16#5C#, 8);
  gmul3_13(52) <= to_unsigned(16#5F#, 8);
  gmul3_13(53) <= to_unsigned(16#5A#, 8);
  gmul3_13(54) <= to_unsigned(16#59#, 8);
  gmul3_13(55) <= to_unsigned(16#48#, 8);
  gmul3_13(56) <= to_unsigned(16#4B#, 8);
  gmul3_13(57) <= to_unsigned(16#4E#, 8);
  gmul3_13(58) <= to_unsigned(16#4D#, 8);
  gmul3_13(59) <= to_unsigned(16#44#, 8);
  gmul3_13(60) <= to_unsigned(16#47#, 8);
  gmul3_13(61) <= to_unsigned(16#42#, 8);
  gmul3_13(62) <= to_unsigned(16#41#, 8);
  gmul3_13(63) <= to_unsigned(16#C0#, 8);
  gmul3_13(64) <= to_unsigned(16#C3#, 8);
  gmul3_13(65) <= to_unsigned(16#C6#, 8);
  gmul3_13(66) <= to_unsigned(16#C5#, 8);
  gmul3_13(67) <= to_unsigned(16#CC#, 8);
  gmul3_13(68) <= to_unsigned(16#CF#, 8);
  gmul3_13(69) <= to_unsigned(16#CA#, 8);
  gmul3_13(70) <= to_unsigned(16#C9#, 8);
  gmul3_13(71) <= to_unsigned(16#D8#, 8);
  gmul3_13(72) <= to_unsigned(16#DB#, 8);
  gmul3_13(73) <= to_unsigned(16#DE#, 8);
  gmul3_13(74) <= to_unsigned(16#DD#, 8);
  gmul3_13(75) <= to_unsigned(16#D4#, 8);
  gmul3_13(76) <= to_unsigned(16#D7#, 8);
  gmul3_13(77) <= to_unsigned(16#D2#, 8);
  gmul3_13(78) <= to_unsigned(16#D1#, 8);
  gmul3_13(79) <= to_unsigned(16#F0#, 8);
  gmul3_13(80) <= to_unsigned(16#F3#, 8);
  gmul3_13(81) <= to_unsigned(16#F6#, 8);
  gmul3_13(82) <= to_unsigned(16#F5#, 8);
  gmul3_13(83) <= to_unsigned(16#FC#, 8);
  gmul3_13(84) <= to_unsigned(16#FF#, 8);
  gmul3_13(85) <= to_unsigned(16#FA#, 8);
  gmul3_13(86) <= to_unsigned(16#F9#, 8);
  gmul3_13(87) <= to_unsigned(16#E8#, 8);
  gmul3_13(88) <= to_unsigned(16#EB#, 8);
  gmul3_13(89) <= to_unsigned(16#EE#, 8);
  gmul3_13(90) <= to_unsigned(16#ED#, 8);
  gmul3_13(91) <= to_unsigned(16#E4#, 8);
  gmul3_13(92) <= to_unsigned(16#E7#, 8);
  gmul3_13(93) <= to_unsigned(16#E2#, 8);
  gmul3_13(94) <= to_unsigned(16#E1#, 8);
  gmul3_13(95) <= to_unsigned(16#A0#, 8);
  gmul3_13(96) <= to_unsigned(16#A3#, 8);
  gmul3_13(97) <= to_unsigned(16#A6#, 8);
  gmul3_13(98) <= to_unsigned(16#A5#, 8);
  gmul3_13(99) <= to_unsigned(16#AC#, 8);
  gmul3_13(100) <= to_unsigned(16#AF#, 8);
  gmul3_13(101) <= to_unsigned(16#AA#, 8);
  gmul3_13(102) <= to_unsigned(16#A9#, 8);
  gmul3_13(103) <= to_unsigned(16#B8#, 8);
  gmul3_13(104) <= to_unsigned(16#BB#, 8);
  gmul3_13(105) <= to_unsigned(16#BE#, 8);
  gmul3_13(106) <= to_unsigned(16#BD#, 8);
  gmul3_13(107) <= to_unsigned(16#B4#, 8);
  gmul3_13(108) <= to_unsigned(16#B7#, 8);
  gmul3_13(109) <= to_unsigned(16#B2#, 8);
  gmul3_13(110) <= to_unsigned(16#B1#, 8);
  gmul3_13(111) <= to_unsigned(16#90#, 8);
  gmul3_13(112) <= to_unsigned(16#93#, 8);
  gmul3_13(113) <= to_unsigned(16#96#, 8);
  gmul3_13(114) <= to_unsigned(16#95#, 8);
  gmul3_13(115) <= to_unsigned(16#9C#, 8);
  gmul3_13(116) <= to_unsigned(16#9F#, 8);
  gmul3_13(117) <= to_unsigned(16#9A#, 8);
  gmul3_13(118) <= to_unsigned(16#99#, 8);
  gmul3_13(119) <= to_unsigned(16#88#, 8);
  gmul3_13(120) <= to_unsigned(16#8B#, 8);
  gmul3_13(121) <= to_unsigned(16#8E#, 8);
  gmul3_13(122) <= to_unsigned(16#8D#, 8);
  gmul3_13(123) <= to_unsigned(16#84#, 8);
  gmul3_13(124) <= to_unsigned(16#87#, 8);
  gmul3_13(125) <= to_unsigned(16#82#, 8);
  gmul3_13(126) <= to_unsigned(16#81#, 8);
  gmul3_13(127) <= to_unsigned(16#9B#, 8);
  gmul3_13(128) <= to_unsigned(16#98#, 8);
  gmul3_13(129) <= to_unsigned(16#9D#, 8);
  gmul3_13(130) <= to_unsigned(16#9E#, 8);
  gmul3_13(131) <= to_unsigned(16#97#, 8);
  gmul3_13(132) <= to_unsigned(16#94#, 8);
  gmul3_13(133) <= to_unsigned(16#91#, 8);
  gmul3_13(134) <= to_unsigned(16#92#, 8);
  gmul3_13(135) <= to_unsigned(16#83#, 8);
  gmul3_13(136) <= to_unsigned(16#80#, 8);
  gmul3_13(137) <= to_unsigned(16#85#, 8);
  gmul3_13(138) <= to_unsigned(16#86#, 8);
  gmul3_13(139) <= to_unsigned(16#8F#, 8);
  gmul3_13(140) <= to_unsigned(16#8C#, 8);
  gmul3_13(141) <= to_unsigned(16#89#, 8);
  gmul3_13(142) <= to_unsigned(16#8A#, 8);
  gmul3_13(143) <= to_unsigned(16#AB#, 8);
  gmul3_13(144) <= to_unsigned(16#A8#, 8);
  gmul3_13(145) <= to_unsigned(16#AD#, 8);
  gmul3_13(146) <= to_unsigned(16#AE#, 8);
  gmul3_13(147) <= to_unsigned(16#A7#, 8);
  gmul3_13(148) <= to_unsigned(16#A4#, 8);
  gmul3_13(149) <= to_unsigned(16#A1#, 8);
  gmul3_13(150) <= to_unsigned(16#A2#, 8);
  gmul3_13(151) <= to_unsigned(16#B3#, 8);
  gmul3_13(152) <= to_unsigned(16#B0#, 8);
  gmul3_13(153) <= to_unsigned(16#B5#, 8);
  gmul3_13(154) <= to_unsigned(16#B6#, 8);
  gmul3_13(155) <= to_unsigned(16#BF#, 8);
  gmul3_13(156) <= to_unsigned(16#BC#, 8);
  gmul3_13(157) <= to_unsigned(16#B9#, 8);
  gmul3_13(158) <= to_unsigned(16#BA#, 8);
  gmul3_13(159) <= to_unsigned(16#FB#, 8);
  gmul3_13(160) <= to_unsigned(16#F8#, 8);
  gmul3_13(161) <= to_unsigned(16#FD#, 8);
  gmul3_13(162) <= to_unsigned(16#FE#, 8);
  gmul3_13(163) <= to_unsigned(16#F7#, 8);
  gmul3_13(164) <= to_unsigned(16#F4#, 8);
  gmul3_13(165) <= to_unsigned(16#F1#, 8);
  gmul3_13(166) <= to_unsigned(16#F2#, 8);
  gmul3_13(167) <= to_unsigned(16#E3#, 8);
  gmul3_13(168) <= to_unsigned(16#E0#, 8);
  gmul3_13(169) <= to_unsigned(16#E5#, 8);
  gmul3_13(170) <= to_unsigned(16#E6#, 8);
  gmul3_13(171) <= to_unsigned(16#EF#, 8);
  gmul3_13(172) <= to_unsigned(16#EC#, 8);
  gmul3_13(173) <= to_unsigned(16#E9#, 8);
  gmul3_13(174) <= to_unsigned(16#EA#, 8);
  gmul3_13(175) <= to_unsigned(16#CB#, 8);
  gmul3_13(176) <= to_unsigned(16#C8#, 8);
  gmul3_13(177) <= to_unsigned(16#CD#, 8);
  gmul3_13(178) <= to_unsigned(16#CE#, 8);
  gmul3_13(179) <= to_unsigned(16#C7#, 8);
  gmul3_13(180) <= to_unsigned(16#C4#, 8);
  gmul3_13(181) <= to_unsigned(16#C1#, 8);
  gmul3_13(182) <= to_unsigned(16#C2#, 8);
  gmul3_13(183) <= to_unsigned(16#D3#, 8);
  gmul3_13(184) <= to_unsigned(16#D0#, 8);
  gmul3_13(185) <= to_unsigned(16#D5#, 8);
  gmul3_13(186) <= to_unsigned(16#D6#, 8);
  gmul3_13(187) <= to_unsigned(16#DF#, 8);
  gmul3_13(188) <= to_unsigned(16#DC#, 8);
  gmul3_13(189) <= to_unsigned(16#D9#, 8);
  gmul3_13(190) <= to_unsigned(16#DA#, 8);
  gmul3_13(191) <= to_unsigned(16#5B#, 8);
  gmul3_13(192) <= to_unsigned(16#58#, 8);
  gmul3_13(193) <= to_unsigned(16#5D#, 8);
  gmul3_13(194) <= to_unsigned(16#5E#, 8);
  gmul3_13(195) <= to_unsigned(16#57#, 8);
  gmul3_13(196) <= to_unsigned(16#54#, 8);
  gmul3_13(197) <= to_unsigned(16#51#, 8);
  gmul3_13(198) <= to_unsigned(16#52#, 8);
  gmul3_13(199) <= to_unsigned(16#43#, 8);
  gmul3_13(200) <= to_unsigned(16#40#, 8);
  gmul3_13(201) <= to_unsigned(16#45#, 8);
  gmul3_13(202) <= to_unsigned(16#46#, 8);
  gmul3_13(203) <= to_unsigned(16#4F#, 8);
  gmul3_13(204) <= to_unsigned(16#4C#, 8);
  gmul3_13(205) <= to_unsigned(16#49#, 8);
  gmul3_13(206) <= to_unsigned(16#4A#, 8);
  gmul3_13(207) <= to_unsigned(16#6B#, 8);
  gmul3_13(208) <= to_unsigned(16#68#, 8);
  gmul3_13(209) <= to_unsigned(16#6D#, 8);
  gmul3_13(210) <= to_unsigned(16#6E#, 8);
  gmul3_13(211) <= to_unsigned(16#67#, 8);
  gmul3_13(212) <= to_unsigned(16#64#, 8);
  gmul3_13(213) <= to_unsigned(16#61#, 8);
  gmul3_13(214) <= to_unsigned(16#62#, 8);
  gmul3_13(215) <= to_unsigned(16#73#, 8);
  gmul3_13(216) <= to_unsigned(16#70#, 8);
  gmul3_13(217) <= to_unsigned(16#75#, 8);
  gmul3_13(218) <= to_unsigned(16#76#, 8);
  gmul3_13(219) <= to_unsigned(16#7F#, 8);
  gmul3_13(220) <= to_unsigned(16#7C#, 8);
  gmul3_13(221) <= to_unsigned(16#79#, 8);
  gmul3_13(222) <= to_unsigned(16#7A#, 8);
  gmul3_13(223) <= to_unsigned(16#3B#, 8);
  gmul3_13(224) <= to_unsigned(16#38#, 8);
  gmul3_13(225) <= to_unsigned(16#3D#, 8);
  gmul3_13(226) <= to_unsigned(16#3E#, 8);
  gmul3_13(227) <= to_unsigned(16#37#, 8);
  gmul3_13(228) <= to_unsigned(16#34#, 8);
  gmul3_13(229) <= to_unsigned(16#31#, 8);
  gmul3_13(230) <= to_unsigned(16#32#, 8);
  gmul3_13(231) <= to_unsigned(16#23#, 8);
  gmul3_13(232) <= to_unsigned(16#20#, 8);
  gmul3_13(233) <= to_unsigned(16#25#, 8);
  gmul3_13(234) <= to_unsigned(16#26#, 8);
  gmul3_13(235) <= to_unsigned(16#2F#, 8);
  gmul3_13(236) <= to_unsigned(16#2C#, 8);
  gmul3_13(237) <= to_unsigned(16#29#, 8);
  gmul3_13(238) <= to_unsigned(16#2A#, 8);
  gmul3_13(239) <= to_unsigned(16#0B#, 8);
  gmul3_13(240) <= to_unsigned(16#08#, 8);
  gmul3_13(241) <= to_unsigned(16#0D#, 8);
  gmul3_13(242) <= to_unsigned(16#0E#, 8);
  gmul3_13(243) <= to_unsigned(16#07#, 8);
  gmul3_13(244) <= to_unsigned(16#04#, 8);
  gmul3_13(245) <= to_unsigned(16#01#, 8);
  gmul3_13(246) <= to_unsigned(16#02#, 8);
  gmul3_13(247) <= to_unsigned(16#13#, 8);
  gmul3_13(248) <= to_unsigned(16#10#, 8);
  gmul3_13(249) <= to_unsigned(16#15#, 8);
  gmul3_13(250) <= to_unsigned(16#16#, 8);
  gmul3_13(251) <= to_unsigned(16#1F#, 8);
  gmul3_13(252) <= to_unsigned(16#1C#, 8);
  gmul3_13(253) <= to_unsigned(16#19#, 8);
  gmul3_13(254) <= to_unsigned(16#1A#, 8);
  gmul3_13(255) <= to_unsigned(16#1A#, 8);

  gmul2_14(0) <= to_unsigned(16#02#, 8);
  gmul2_14(1) <= to_unsigned(16#04#, 8);
  gmul2_14(2) <= to_unsigned(16#06#, 8);
  gmul2_14(3) <= to_unsigned(16#08#, 8);
  gmul2_14(4) <= to_unsigned(16#0A#, 8);
  gmul2_14(5) <= to_unsigned(16#0C#, 8);
  gmul2_14(6) <= to_unsigned(16#0E#, 8);
  gmul2_14(7) <= to_unsigned(16#10#, 8);
  gmul2_14(8) <= to_unsigned(16#12#, 8);
  gmul2_14(9) <= to_unsigned(16#14#, 8);
  gmul2_14(10) <= to_unsigned(16#16#, 8);
  gmul2_14(11) <= to_unsigned(16#18#, 8);
  gmul2_14(12) <= to_unsigned(16#1A#, 8);
  gmul2_14(13) <= to_unsigned(16#1C#, 8);
  gmul2_14(14) <= to_unsigned(16#1E#, 8);
  gmul2_14(15) <= to_unsigned(16#20#, 8);
  gmul2_14(16) <= to_unsigned(16#22#, 8);
  gmul2_14(17) <= to_unsigned(16#24#, 8);
  gmul2_14(18) <= to_unsigned(16#26#, 8);
  gmul2_14(19) <= to_unsigned(16#28#, 8);
  gmul2_14(20) <= to_unsigned(16#2A#, 8);
  gmul2_14(21) <= to_unsigned(16#2C#, 8);
  gmul2_14(22) <= to_unsigned(16#2E#, 8);
  gmul2_14(23) <= to_unsigned(16#30#, 8);
  gmul2_14(24) <= to_unsigned(16#32#, 8);
  gmul2_14(25) <= to_unsigned(16#34#, 8);
  gmul2_14(26) <= to_unsigned(16#36#, 8);
  gmul2_14(27) <= to_unsigned(16#38#, 8);
  gmul2_14(28) <= to_unsigned(16#3A#, 8);
  gmul2_14(29) <= to_unsigned(16#3C#, 8);
  gmul2_14(30) <= to_unsigned(16#3E#, 8);
  gmul2_14(31) <= to_unsigned(16#40#, 8);
  gmul2_14(32) <= to_unsigned(16#42#, 8);
  gmul2_14(33) <= to_unsigned(16#44#, 8);
  gmul2_14(34) <= to_unsigned(16#46#, 8);
  gmul2_14(35) <= to_unsigned(16#48#, 8);
  gmul2_14(36) <= to_unsigned(16#4A#, 8);
  gmul2_14(37) <= to_unsigned(16#4C#, 8);
  gmul2_14(38) <= to_unsigned(16#4E#, 8);
  gmul2_14(39) <= to_unsigned(16#50#, 8);
  gmul2_14(40) <= to_unsigned(16#52#, 8);
  gmul2_14(41) <= to_unsigned(16#54#, 8);
  gmul2_14(42) <= to_unsigned(16#56#, 8);
  gmul2_14(43) <= to_unsigned(16#58#, 8);
  gmul2_14(44) <= to_unsigned(16#5A#, 8);
  gmul2_14(45) <= to_unsigned(16#5C#, 8);
  gmul2_14(46) <= to_unsigned(16#5E#, 8);
  gmul2_14(47) <= to_unsigned(16#60#, 8);
  gmul2_14(48) <= to_unsigned(16#62#, 8);
  gmul2_14(49) <= to_unsigned(16#64#, 8);
  gmul2_14(50) <= to_unsigned(16#66#, 8);
  gmul2_14(51) <= to_unsigned(16#68#, 8);
  gmul2_14(52) <= to_unsigned(16#6A#, 8);
  gmul2_14(53) <= to_unsigned(16#6C#, 8);
  gmul2_14(54) <= to_unsigned(16#6E#, 8);
  gmul2_14(55) <= to_unsigned(16#70#, 8);
  gmul2_14(56) <= to_unsigned(16#72#, 8);
  gmul2_14(57) <= to_unsigned(16#74#, 8);
  gmul2_14(58) <= to_unsigned(16#76#, 8);
  gmul2_14(59) <= to_unsigned(16#78#, 8);
  gmul2_14(60) <= to_unsigned(16#7A#, 8);
  gmul2_14(61) <= to_unsigned(16#7C#, 8);
  gmul2_14(62) <= to_unsigned(16#7E#, 8);
  gmul2_14(63) <= to_unsigned(16#80#, 8);
  gmul2_14(64) <= to_unsigned(16#82#, 8);
  gmul2_14(65) <= to_unsigned(16#84#, 8);
  gmul2_14(66) <= to_unsigned(16#86#, 8);
  gmul2_14(67) <= to_unsigned(16#88#, 8);
  gmul2_14(68) <= to_unsigned(16#8A#, 8);
  gmul2_14(69) <= to_unsigned(16#8C#, 8);
  gmul2_14(70) <= to_unsigned(16#8E#, 8);
  gmul2_14(71) <= to_unsigned(16#90#, 8);
  gmul2_14(72) <= to_unsigned(16#92#, 8);
  gmul2_14(73) <= to_unsigned(16#94#, 8);
  gmul2_14(74) <= to_unsigned(16#96#, 8);
  gmul2_14(75) <= to_unsigned(16#98#, 8);
  gmul2_14(76) <= to_unsigned(16#9A#, 8);
  gmul2_14(77) <= to_unsigned(16#9C#, 8);
  gmul2_14(78) <= to_unsigned(16#9E#, 8);
  gmul2_14(79) <= to_unsigned(16#A0#, 8);
  gmul2_14(80) <= to_unsigned(16#A2#, 8);
  gmul2_14(81) <= to_unsigned(16#A4#, 8);
  gmul2_14(82) <= to_unsigned(16#A6#, 8);
  gmul2_14(83) <= to_unsigned(16#A8#, 8);
  gmul2_14(84) <= to_unsigned(16#AA#, 8);
  gmul2_14(85) <= to_unsigned(16#AC#, 8);
  gmul2_14(86) <= to_unsigned(16#AE#, 8);
  gmul2_14(87) <= to_unsigned(16#B0#, 8);
  gmul2_14(88) <= to_unsigned(16#B2#, 8);
  gmul2_14(89) <= to_unsigned(16#B4#, 8);
  gmul2_14(90) <= to_unsigned(16#B6#, 8);
  gmul2_14(91) <= to_unsigned(16#B8#, 8);
  gmul2_14(92) <= to_unsigned(16#BA#, 8);
  gmul2_14(93) <= to_unsigned(16#BC#, 8);
  gmul2_14(94) <= to_unsigned(16#BE#, 8);
  gmul2_14(95) <= to_unsigned(16#C0#, 8);
  gmul2_14(96) <= to_unsigned(16#C2#, 8);
  gmul2_14(97) <= to_unsigned(16#C4#, 8);
  gmul2_14(98) <= to_unsigned(16#C6#, 8);
  gmul2_14(99) <= to_unsigned(16#C8#, 8);
  gmul2_14(100) <= to_unsigned(16#CA#, 8);
  gmul2_14(101) <= to_unsigned(16#CC#, 8);
  gmul2_14(102) <= to_unsigned(16#CE#, 8);
  gmul2_14(103) <= to_unsigned(16#D0#, 8);
  gmul2_14(104) <= to_unsigned(16#D2#, 8);
  gmul2_14(105) <= to_unsigned(16#D4#, 8);
  gmul2_14(106) <= to_unsigned(16#D6#, 8);
  gmul2_14(107) <= to_unsigned(16#D8#, 8);
  gmul2_14(108) <= to_unsigned(16#DA#, 8);
  gmul2_14(109) <= to_unsigned(16#DC#, 8);
  gmul2_14(110) <= to_unsigned(16#DE#, 8);
  gmul2_14(111) <= to_unsigned(16#E0#, 8);
  gmul2_14(112) <= to_unsigned(16#E2#, 8);
  gmul2_14(113) <= to_unsigned(16#E4#, 8);
  gmul2_14(114) <= to_unsigned(16#E6#, 8);
  gmul2_14(115) <= to_unsigned(16#E8#, 8);
  gmul2_14(116) <= to_unsigned(16#EA#, 8);
  gmul2_14(117) <= to_unsigned(16#EC#, 8);
  gmul2_14(118) <= to_unsigned(16#EE#, 8);
  gmul2_14(119) <= to_unsigned(16#F0#, 8);
  gmul2_14(120) <= to_unsigned(16#F2#, 8);
  gmul2_14(121) <= to_unsigned(16#F4#, 8);
  gmul2_14(122) <= to_unsigned(16#F6#, 8);
  gmul2_14(123) <= to_unsigned(16#F8#, 8);
  gmul2_14(124) <= to_unsigned(16#FA#, 8);
  gmul2_14(125) <= to_unsigned(16#FC#, 8);
  gmul2_14(126) <= to_unsigned(16#FE#, 8);
  gmul2_14(127) <= to_unsigned(16#1B#, 8);
  gmul2_14(128) <= to_unsigned(16#19#, 8);
  gmul2_14(129) <= to_unsigned(16#1F#, 8);
  gmul2_14(130) <= to_unsigned(16#1D#, 8);
  gmul2_14(131) <= to_unsigned(16#13#, 8);
  gmul2_14(132) <= to_unsigned(16#11#, 8);
  gmul2_14(133) <= to_unsigned(16#17#, 8);
  gmul2_14(134) <= to_unsigned(16#15#, 8);
  gmul2_14(135) <= to_unsigned(16#0B#, 8);
  gmul2_14(136) <= to_unsigned(16#09#, 8);
  gmul2_14(137) <= to_unsigned(16#0F#, 8);
  gmul2_14(138) <= to_unsigned(16#0D#, 8);
  gmul2_14(139) <= to_unsigned(16#03#, 8);
  gmul2_14(140) <= to_unsigned(16#01#, 8);
  gmul2_14(141) <= to_unsigned(16#07#, 8);
  gmul2_14(142) <= to_unsigned(16#05#, 8);
  gmul2_14(143) <= to_unsigned(16#3B#, 8);
  gmul2_14(144) <= to_unsigned(16#39#, 8);
  gmul2_14(145) <= to_unsigned(16#3F#, 8);
  gmul2_14(146) <= to_unsigned(16#3D#, 8);
  gmul2_14(147) <= to_unsigned(16#33#, 8);
  gmul2_14(148) <= to_unsigned(16#31#, 8);
  gmul2_14(149) <= to_unsigned(16#37#, 8);
  gmul2_14(150) <= to_unsigned(16#35#, 8);
  gmul2_14(151) <= to_unsigned(16#2B#, 8);
  gmul2_14(152) <= to_unsigned(16#29#, 8);
  gmul2_14(153) <= to_unsigned(16#2F#, 8);
  gmul2_14(154) <= to_unsigned(16#2D#, 8);
  gmul2_14(155) <= to_unsigned(16#23#, 8);
  gmul2_14(156) <= to_unsigned(16#21#, 8);
  gmul2_14(157) <= to_unsigned(16#27#, 8);
  gmul2_14(158) <= to_unsigned(16#25#, 8);
  gmul2_14(159) <= to_unsigned(16#5B#, 8);
  gmul2_14(160) <= to_unsigned(16#59#, 8);
  gmul2_14(161) <= to_unsigned(16#5F#, 8);
  gmul2_14(162) <= to_unsigned(16#5D#, 8);
  gmul2_14(163) <= to_unsigned(16#53#, 8);
  gmul2_14(164) <= to_unsigned(16#51#, 8);
  gmul2_14(165) <= to_unsigned(16#57#, 8);
  gmul2_14(166) <= to_unsigned(16#55#, 8);
  gmul2_14(167) <= to_unsigned(16#4B#, 8);
  gmul2_14(168) <= to_unsigned(16#49#, 8);
  gmul2_14(169) <= to_unsigned(16#4F#, 8);
  gmul2_14(170) <= to_unsigned(16#4D#, 8);
  gmul2_14(171) <= to_unsigned(16#43#, 8);
  gmul2_14(172) <= to_unsigned(16#41#, 8);
  gmul2_14(173) <= to_unsigned(16#47#, 8);
  gmul2_14(174) <= to_unsigned(16#45#, 8);
  gmul2_14(175) <= to_unsigned(16#7B#, 8);
  gmul2_14(176) <= to_unsigned(16#79#, 8);
  gmul2_14(177) <= to_unsigned(16#7F#, 8);
  gmul2_14(178) <= to_unsigned(16#7D#, 8);
  gmul2_14(179) <= to_unsigned(16#73#, 8);
  gmul2_14(180) <= to_unsigned(16#71#, 8);
  gmul2_14(181) <= to_unsigned(16#77#, 8);
  gmul2_14(182) <= to_unsigned(16#75#, 8);
  gmul2_14(183) <= to_unsigned(16#6B#, 8);
  gmul2_14(184) <= to_unsigned(16#69#, 8);
  gmul2_14(185) <= to_unsigned(16#6F#, 8);
  gmul2_14(186) <= to_unsigned(16#6D#, 8);
  gmul2_14(187) <= to_unsigned(16#63#, 8);
  gmul2_14(188) <= to_unsigned(16#61#, 8);
  gmul2_14(189) <= to_unsigned(16#67#, 8);
  gmul2_14(190) <= to_unsigned(16#65#, 8);
  gmul2_14(191) <= to_unsigned(16#9B#, 8);
  gmul2_14(192) <= to_unsigned(16#99#, 8);
  gmul2_14(193) <= to_unsigned(16#9F#, 8);
  gmul2_14(194) <= to_unsigned(16#9D#, 8);
  gmul2_14(195) <= to_unsigned(16#93#, 8);
  gmul2_14(196) <= to_unsigned(16#91#, 8);
  gmul2_14(197) <= to_unsigned(16#97#, 8);
  gmul2_14(198) <= to_unsigned(16#95#, 8);
  gmul2_14(199) <= to_unsigned(16#8B#, 8);
  gmul2_14(200) <= to_unsigned(16#89#, 8);
  gmul2_14(201) <= to_unsigned(16#8F#, 8);
  gmul2_14(202) <= to_unsigned(16#8D#, 8);
  gmul2_14(203) <= to_unsigned(16#83#, 8);
  gmul2_14(204) <= to_unsigned(16#81#, 8);
  gmul2_14(205) <= to_unsigned(16#87#, 8);
  gmul2_14(206) <= to_unsigned(16#85#, 8);
  gmul2_14(207) <= to_unsigned(16#BB#, 8);
  gmul2_14(208) <= to_unsigned(16#B9#, 8);
  gmul2_14(209) <= to_unsigned(16#BF#, 8);
  gmul2_14(210) <= to_unsigned(16#BD#, 8);
  gmul2_14(211) <= to_unsigned(16#B3#, 8);
  gmul2_14(212) <= to_unsigned(16#B1#, 8);
  gmul2_14(213) <= to_unsigned(16#B7#, 8);
  gmul2_14(214) <= to_unsigned(16#B5#, 8);
  gmul2_14(215) <= to_unsigned(16#AB#, 8);
  gmul2_14(216) <= to_unsigned(16#A9#, 8);
  gmul2_14(217) <= to_unsigned(16#AF#, 8);
  gmul2_14(218) <= to_unsigned(16#AD#, 8);
  gmul2_14(219) <= to_unsigned(16#A3#, 8);
  gmul2_14(220) <= to_unsigned(16#A1#, 8);
  gmul2_14(221) <= to_unsigned(16#A7#, 8);
  gmul2_14(222) <= to_unsigned(16#A5#, 8);
  gmul2_14(223) <= to_unsigned(16#DB#, 8);
  gmul2_14(224) <= to_unsigned(16#D9#, 8);
  gmul2_14(225) <= to_unsigned(16#DF#, 8);
  gmul2_14(226) <= to_unsigned(16#DD#, 8);
  gmul2_14(227) <= to_unsigned(16#D3#, 8);
  gmul2_14(228) <= to_unsigned(16#D1#, 8);
  gmul2_14(229) <= to_unsigned(16#D7#, 8);
  gmul2_14(230) <= to_unsigned(16#D5#, 8);
  gmul2_14(231) <= to_unsigned(16#CB#, 8);
  gmul2_14(232) <= to_unsigned(16#C9#, 8);
  gmul2_14(233) <= to_unsigned(16#CF#, 8);
  gmul2_14(234) <= to_unsigned(16#CD#, 8);
  gmul2_14(235) <= to_unsigned(16#C3#, 8);
  gmul2_14(236) <= to_unsigned(16#C1#, 8);
  gmul2_14(237) <= to_unsigned(16#C7#, 8);
  gmul2_14(238) <= to_unsigned(16#C5#, 8);
  gmul2_14(239) <= to_unsigned(16#FB#, 8);
  gmul2_14(240) <= to_unsigned(16#F9#, 8);
  gmul2_14(241) <= to_unsigned(16#FF#, 8);
  gmul2_14(242) <= to_unsigned(16#FD#, 8);
  gmul2_14(243) <= to_unsigned(16#F3#, 8);
  gmul2_14(244) <= to_unsigned(16#F1#, 8);
  gmul2_14(245) <= to_unsigned(16#F7#, 8);
  gmul2_14(246) <= to_unsigned(16#F5#, 8);
  gmul2_14(247) <= to_unsigned(16#EB#, 8);
  gmul2_14(248) <= to_unsigned(16#E9#, 8);
  gmul2_14(249) <= to_unsigned(16#EF#, 8);
  gmul2_14(250) <= to_unsigned(16#ED#, 8);
  gmul2_14(251) <= to_unsigned(16#E3#, 8);
  gmul2_14(252) <= to_unsigned(16#E1#, 8);
  gmul2_14(253) <= to_unsigned(16#E7#, 8);
  gmul2_14(254) <= to_unsigned(16#E5#, 8);
  gmul2_14(255) <= to_unsigned(16#E5#, 8);

  gmul3_14(0) <= to_unsigned(16#03#, 8);
  gmul3_14(1) <= to_unsigned(16#06#, 8);
  gmul3_14(2) <= to_unsigned(16#05#, 8);
  gmul3_14(3) <= to_unsigned(16#0C#, 8);
  gmul3_14(4) <= to_unsigned(16#0F#, 8);
  gmul3_14(5) <= to_unsigned(16#0A#, 8);
  gmul3_14(6) <= to_unsigned(16#09#, 8);
  gmul3_14(7) <= to_unsigned(16#18#, 8);
  gmul3_14(8) <= to_unsigned(16#1B#, 8);
  gmul3_14(9) <= to_unsigned(16#1E#, 8);
  gmul3_14(10) <= to_unsigned(16#1D#, 8);
  gmul3_14(11) <= to_unsigned(16#14#, 8);
  gmul3_14(12) <= to_unsigned(16#17#, 8);
  gmul3_14(13) <= to_unsigned(16#12#, 8);
  gmul3_14(14) <= to_unsigned(16#11#, 8);
  gmul3_14(15) <= to_unsigned(16#30#, 8);
  gmul3_14(16) <= to_unsigned(16#33#, 8);
  gmul3_14(17) <= to_unsigned(16#36#, 8);
  gmul3_14(18) <= to_unsigned(16#35#, 8);
  gmul3_14(19) <= to_unsigned(16#3C#, 8);
  gmul3_14(20) <= to_unsigned(16#3F#, 8);
  gmul3_14(21) <= to_unsigned(16#3A#, 8);
  gmul3_14(22) <= to_unsigned(16#39#, 8);
  gmul3_14(23) <= to_unsigned(16#28#, 8);
  gmul3_14(24) <= to_unsigned(16#2B#, 8);
  gmul3_14(25) <= to_unsigned(16#2E#, 8);
  gmul3_14(26) <= to_unsigned(16#2D#, 8);
  gmul3_14(27) <= to_unsigned(16#24#, 8);
  gmul3_14(28) <= to_unsigned(16#27#, 8);
  gmul3_14(29) <= to_unsigned(16#22#, 8);
  gmul3_14(30) <= to_unsigned(16#21#, 8);
  gmul3_14(31) <= to_unsigned(16#60#, 8);
  gmul3_14(32) <= to_unsigned(16#63#, 8);
  gmul3_14(33) <= to_unsigned(16#66#, 8);
  gmul3_14(34) <= to_unsigned(16#65#, 8);
  gmul3_14(35) <= to_unsigned(16#6C#, 8);
  gmul3_14(36) <= to_unsigned(16#6F#, 8);
  gmul3_14(37) <= to_unsigned(16#6A#, 8);
  gmul3_14(38) <= to_unsigned(16#69#, 8);
  gmul3_14(39) <= to_unsigned(16#78#, 8);
  gmul3_14(40) <= to_unsigned(16#7B#, 8);
  gmul3_14(41) <= to_unsigned(16#7E#, 8);
  gmul3_14(42) <= to_unsigned(16#7D#, 8);
  gmul3_14(43) <= to_unsigned(16#74#, 8);
  gmul3_14(44) <= to_unsigned(16#77#, 8);
  gmul3_14(45) <= to_unsigned(16#72#, 8);
  gmul3_14(46) <= to_unsigned(16#71#, 8);
  gmul3_14(47) <= to_unsigned(16#50#, 8);
  gmul3_14(48) <= to_unsigned(16#53#, 8);
  gmul3_14(49) <= to_unsigned(16#56#, 8);
  gmul3_14(50) <= to_unsigned(16#55#, 8);
  gmul3_14(51) <= to_unsigned(16#5C#, 8);
  gmul3_14(52) <= to_unsigned(16#5F#, 8);
  gmul3_14(53) <= to_unsigned(16#5A#, 8);
  gmul3_14(54) <= to_unsigned(16#59#, 8);
  gmul3_14(55) <= to_unsigned(16#48#, 8);
  gmul3_14(56) <= to_unsigned(16#4B#, 8);
  gmul3_14(57) <= to_unsigned(16#4E#, 8);
  gmul3_14(58) <= to_unsigned(16#4D#, 8);
  gmul3_14(59) <= to_unsigned(16#44#, 8);
  gmul3_14(60) <= to_unsigned(16#47#, 8);
  gmul3_14(61) <= to_unsigned(16#42#, 8);
  gmul3_14(62) <= to_unsigned(16#41#, 8);
  gmul3_14(63) <= to_unsigned(16#C0#, 8);
  gmul3_14(64) <= to_unsigned(16#C3#, 8);
  gmul3_14(65) <= to_unsigned(16#C6#, 8);
  gmul3_14(66) <= to_unsigned(16#C5#, 8);
  gmul3_14(67) <= to_unsigned(16#CC#, 8);
  gmul3_14(68) <= to_unsigned(16#CF#, 8);
  gmul3_14(69) <= to_unsigned(16#CA#, 8);
  gmul3_14(70) <= to_unsigned(16#C9#, 8);
  gmul3_14(71) <= to_unsigned(16#D8#, 8);
  gmul3_14(72) <= to_unsigned(16#DB#, 8);
  gmul3_14(73) <= to_unsigned(16#DE#, 8);
  gmul3_14(74) <= to_unsigned(16#DD#, 8);
  gmul3_14(75) <= to_unsigned(16#D4#, 8);
  gmul3_14(76) <= to_unsigned(16#D7#, 8);
  gmul3_14(77) <= to_unsigned(16#D2#, 8);
  gmul3_14(78) <= to_unsigned(16#D1#, 8);
  gmul3_14(79) <= to_unsigned(16#F0#, 8);
  gmul3_14(80) <= to_unsigned(16#F3#, 8);
  gmul3_14(81) <= to_unsigned(16#F6#, 8);
  gmul3_14(82) <= to_unsigned(16#F5#, 8);
  gmul3_14(83) <= to_unsigned(16#FC#, 8);
  gmul3_14(84) <= to_unsigned(16#FF#, 8);
  gmul3_14(85) <= to_unsigned(16#FA#, 8);
  gmul3_14(86) <= to_unsigned(16#F9#, 8);
  gmul3_14(87) <= to_unsigned(16#E8#, 8);
  gmul3_14(88) <= to_unsigned(16#EB#, 8);
  gmul3_14(89) <= to_unsigned(16#EE#, 8);
  gmul3_14(90) <= to_unsigned(16#ED#, 8);
  gmul3_14(91) <= to_unsigned(16#E4#, 8);
  gmul3_14(92) <= to_unsigned(16#E7#, 8);
  gmul3_14(93) <= to_unsigned(16#E2#, 8);
  gmul3_14(94) <= to_unsigned(16#E1#, 8);
  gmul3_14(95) <= to_unsigned(16#A0#, 8);
  gmul3_14(96) <= to_unsigned(16#A3#, 8);
  gmul3_14(97) <= to_unsigned(16#A6#, 8);
  gmul3_14(98) <= to_unsigned(16#A5#, 8);
  gmul3_14(99) <= to_unsigned(16#AC#, 8);
  gmul3_14(100) <= to_unsigned(16#AF#, 8);
  gmul3_14(101) <= to_unsigned(16#AA#, 8);
  gmul3_14(102) <= to_unsigned(16#A9#, 8);
  gmul3_14(103) <= to_unsigned(16#B8#, 8);
  gmul3_14(104) <= to_unsigned(16#BB#, 8);
  gmul3_14(105) <= to_unsigned(16#BE#, 8);
  gmul3_14(106) <= to_unsigned(16#BD#, 8);
  gmul3_14(107) <= to_unsigned(16#B4#, 8);
  gmul3_14(108) <= to_unsigned(16#B7#, 8);
  gmul3_14(109) <= to_unsigned(16#B2#, 8);
  gmul3_14(110) <= to_unsigned(16#B1#, 8);
  gmul3_14(111) <= to_unsigned(16#90#, 8);
  gmul3_14(112) <= to_unsigned(16#93#, 8);
  gmul3_14(113) <= to_unsigned(16#96#, 8);
  gmul3_14(114) <= to_unsigned(16#95#, 8);
  gmul3_14(115) <= to_unsigned(16#9C#, 8);
  gmul3_14(116) <= to_unsigned(16#9F#, 8);
  gmul3_14(117) <= to_unsigned(16#9A#, 8);
  gmul3_14(118) <= to_unsigned(16#99#, 8);
  gmul3_14(119) <= to_unsigned(16#88#, 8);
  gmul3_14(120) <= to_unsigned(16#8B#, 8);
  gmul3_14(121) <= to_unsigned(16#8E#, 8);
  gmul3_14(122) <= to_unsigned(16#8D#, 8);
  gmul3_14(123) <= to_unsigned(16#84#, 8);
  gmul3_14(124) <= to_unsigned(16#87#, 8);
  gmul3_14(125) <= to_unsigned(16#82#, 8);
  gmul3_14(126) <= to_unsigned(16#81#, 8);
  gmul3_14(127) <= to_unsigned(16#9B#, 8);
  gmul3_14(128) <= to_unsigned(16#98#, 8);
  gmul3_14(129) <= to_unsigned(16#9D#, 8);
  gmul3_14(130) <= to_unsigned(16#9E#, 8);
  gmul3_14(131) <= to_unsigned(16#97#, 8);
  gmul3_14(132) <= to_unsigned(16#94#, 8);
  gmul3_14(133) <= to_unsigned(16#91#, 8);
  gmul3_14(134) <= to_unsigned(16#92#, 8);
  gmul3_14(135) <= to_unsigned(16#83#, 8);
  gmul3_14(136) <= to_unsigned(16#80#, 8);
  gmul3_14(137) <= to_unsigned(16#85#, 8);
  gmul3_14(138) <= to_unsigned(16#86#, 8);
  gmul3_14(139) <= to_unsigned(16#8F#, 8);
  gmul3_14(140) <= to_unsigned(16#8C#, 8);
  gmul3_14(141) <= to_unsigned(16#89#, 8);
  gmul3_14(142) <= to_unsigned(16#8A#, 8);
  gmul3_14(143) <= to_unsigned(16#AB#, 8);
  gmul3_14(144) <= to_unsigned(16#A8#, 8);
  gmul3_14(145) <= to_unsigned(16#AD#, 8);
  gmul3_14(146) <= to_unsigned(16#AE#, 8);
  gmul3_14(147) <= to_unsigned(16#A7#, 8);
  gmul3_14(148) <= to_unsigned(16#A4#, 8);
  gmul3_14(149) <= to_unsigned(16#A1#, 8);
  gmul3_14(150) <= to_unsigned(16#A2#, 8);
  gmul3_14(151) <= to_unsigned(16#B3#, 8);
  gmul3_14(152) <= to_unsigned(16#B0#, 8);
  gmul3_14(153) <= to_unsigned(16#B5#, 8);
  gmul3_14(154) <= to_unsigned(16#B6#, 8);
  gmul3_14(155) <= to_unsigned(16#BF#, 8);
  gmul3_14(156) <= to_unsigned(16#BC#, 8);
  gmul3_14(157) <= to_unsigned(16#B9#, 8);
  gmul3_14(158) <= to_unsigned(16#BA#, 8);
  gmul3_14(159) <= to_unsigned(16#FB#, 8);
  gmul3_14(160) <= to_unsigned(16#F8#, 8);
  gmul3_14(161) <= to_unsigned(16#FD#, 8);
  gmul3_14(162) <= to_unsigned(16#FE#, 8);
  gmul3_14(163) <= to_unsigned(16#F7#, 8);
  gmul3_14(164) <= to_unsigned(16#F4#, 8);
  gmul3_14(165) <= to_unsigned(16#F1#, 8);
  gmul3_14(166) <= to_unsigned(16#F2#, 8);
  gmul3_14(167) <= to_unsigned(16#E3#, 8);
  gmul3_14(168) <= to_unsigned(16#E0#, 8);
  gmul3_14(169) <= to_unsigned(16#E5#, 8);
  gmul3_14(170) <= to_unsigned(16#E6#, 8);
  gmul3_14(171) <= to_unsigned(16#EF#, 8);
  gmul3_14(172) <= to_unsigned(16#EC#, 8);
  gmul3_14(173) <= to_unsigned(16#E9#, 8);
  gmul3_14(174) <= to_unsigned(16#EA#, 8);
  gmul3_14(175) <= to_unsigned(16#CB#, 8);
  gmul3_14(176) <= to_unsigned(16#C8#, 8);
  gmul3_14(177) <= to_unsigned(16#CD#, 8);
  gmul3_14(178) <= to_unsigned(16#CE#, 8);
  gmul3_14(179) <= to_unsigned(16#C7#, 8);
  gmul3_14(180) <= to_unsigned(16#C4#, 8);
  gmul3_14(181) <= to_unsigned(16#C1#, 8);
  gmul3_14(182) <= to_unsigned(16#C2#, 8);
  gmul3_14(183) <= to_unsigned(16#D3#, 8);
  gmul3_14(184) <= to_unsigned(16#D0#, 8);
  gmul3_14(185) <= to_unsigned(16#D5#, 8);
  gmul3_14(186) <= to_unsigned(16#D6#, 8);
  gmul3_14(187) <= to_unsigned(16#DF#, 8);
  gmul3_14(188) <= to_unsigned(16#DC#, 8);
  gmul3_14(189) <= to_unsigned(16#D9#, 8);
  gmul3_14(190) <= to_unsigned(16#DA#, 8);
  gmul3_14(191) <= to_unsigned(16#5B#, 8);
  gmul3_14(192) <= to_unsigned(16#58#, 8);
  gmul3_14(193) <= to_unsigned(16#5D#, 8);
  gmul3_14(194) <= to_unsigned(16#5E#, 8);
  gmul3_14(195) <= to_unsigned(16#57#, 8);
  gmul3_14(196) <= to_unsigned(16#54#, 8);
  gmul3_14(197) <= to_unsigned(16#51#, 8);
  gmul3_14(198) <= to_unsigned(16#52#, 8);
  gmul3_14(199) <= to_unsigned(16#43#, 8);
  gmul3_14(200) <= to_unsigned(16#40#, 8);
  gmul3_14(201) <= to_unsigned(16#45#, 8);
  gmul3_14(202) <= to_unsigned(16#46#, 8);
  gmul3_14(203) <= to_unsigned(16#4F#, 8);
  gmul3_14(204) <= to_unsigned(16#4C#, 8);
  gmul3_14(205) <= to_unsigned(16#49#, 8);
  gmul3_14(206) <= to_unsigned(16#4A#, 8);
  gmul3_14(207) <= to_unsigned(16#6B#, 8);
  gmul3_14(208) <= to_unsigned(16#68#, 8);
  gmul3_14(209) <= to_unsigned(16#6D#, 8);
  gmul3_14(210) <= to_unsigned(16#6E#, 8);
  gmul3_14(211) <= to_unsigned(16#67#, 8);
  gmul3_14(212) <= to_unsigned(16#64#, 8);
  gmul3_14(213) <= to_unsigned(16#61#, 8);
  gmul3_14(214) <= to_unsigned(16#62#, 8);
  gmul3_14(215) <= to_unsigned(16#73#, 8);
  gmul3_14(216) <= to_unsigned(16#70#, 8);
  gmul3_14(217) <= to_unsigned(16#75#, 8);
  gmul3_14(218) <= to_unsigned(16#76#, 8);
  gmul3_14(219) <= to_unsigned(16#7F#, 8);
  gmul3_14(220) <= to_unsigned(16#7C#, 8);
  gmul3_14(221) <= to_unsigned(16#79#, 8);
  gmul3_14(222) <= to_unsigned(16#7A#, 8);
  gmul3_14(223) <= to_unsigned(16#3B#, 8);
  gmul3_14(224) <= to_unsigned(16#38#, 8);
  gmul3_14(225) <= to_unsigned(16#3D#, 8);
  gmul3_14(226) <= to_unsigned(16#3E#, 8);
  gmul3_14(227) <= to_unsigned(16#37#, 8);
  gmul3_14(228) <= to_unsigned(16#34#, 8);
  gmul3_14(229) <= to_unsigned(16#31#, 8);
  gmul3_14(230) <= to_unsigned(16#32#, 8);
  gmul3_14(231) <= to_unsigned(16#23#, 8);
  gmul3_14(232) <= to_unsigned(16#20#, 8);
  gmul3_14(233) <= to_unsigned(16#25#, 8);
  gmul3_14(234) <= to_unsigned(16#26#, 8);
  gmul3_14(235) <= to_unsigned(16#2F#, 8);
  gmul3_14(236) <= to_unsigned(16#2C#, 8);
  gmul3_14(237) <= to_unsigned(16#29#, 8);
  gmul3_14(238) <= to_unsigned(16#2A#, 8);
  gmul3_14(239) <= to_unsigned(16#0B#, 8);
  gmul3_14(240) <= to_unsigned(16#08#, 8);
  gmul3_14(241) <= to_unsigned(16#0D#, 8);
  gmul3_14(242) <= to_unsigned(16#0E#, 8);
  gmul3_14(243) <= to_unsigned(16#07#, 8);
  gmul3_14(244) <= to_unsigned(16#04#, 8);
  gmul3_14(245) <= to_unsigned(16#01#, 8);
  gmul3_14(246) <= to_unsigned(16#02#, 8);
  gmul3_14(247) <= to_unsigned(16#13#, 8);
  gmul3_14(248) <= to_unsigned(16#10#, 8);
  gmul3_14(249) <= to_unsigned(16#15#, 8);
  gmul3_14(250) <= to_unsigned(16#16#, 8);
  gmul3_14(251) <= to_unsigned(16#1F#, 8);
  gmul3_14(252) <= to_unsigned(16#1C#, 8);
  gmul3_14(253) <= to_unsigned(16#19#, 8);
  gmul3_14(254) <= to_unsigned(16#1A#, 8);
  gmul3_14(255) <= to_unsigned(16#1A#, 8);

  gmul3_15(0) <= to_unsigned(16#03#, 8);
  gmul3_15(1) <= to_unsigned(16#06#, 8);
  gmul3_15(2) <= to_unsigned(16#05#, 8);
  gmul3_15(3) <= to_unsigned(16#0C#, 8);
  gmul3_15(4) <= to_unsigned(16#0F#, 8);
  gmul3_15(5) <= to_unsigned(16#0A#, 8);
  gmul3_15(6) <= to_unsigned(16#09#, 8);
  gmul3_15(7) <= to_unsigned(16#18#, 8);
  gmul3_15(8) <= to_unsigned(16#1B#, 8);
  gmul3_15(9) <= to_unsigned(16#1E#, 8);
  gmul3_15(10) <= to_unsigned(16#1D#, 8);
  gmul3_15(11) <= to_unsigned(16#14#, 8);
  gmul3_15(12) <= to_unsigned(16#17#, 8);
  gmul3_15(13) <= to_unsigned(16#12#, 8);
  gmul3_15(14) <= to_unsigned(16#11#, 8);
  gmul3_15(15) <= to_unsigned(16#30#, 8);
  gmul3_15(16) <= to_unsigned(16#33#, 8);
  gmul3_15(17) <= to_unsigned(16#36#, 8);
  gmul3_15(18) <= to_unsigned(16#35#, 8);
  gmul3_15(19) <= to_unsigned(16#3C#, 8);
  gmul3_15(20) <= to_unsigned(16#3F#, 8);
  gmul3_15(21) <= to_unsigned(16#3A#, 8);
  gmul3_15(22) <= to_unsigned(16#39#, 8);
  gmul3_15(23) <= to_unsigned(16#28#, 8);
  gmul3_15(24) <= to_unsigned(16#2B#, 8);
  gmul3_15(25) <= to_unsigned(16#2E#, 8);
  gmul3_15(26) <= to_unsigned(16#2D#, 8);
  gmul3_15(27) <= to_unsigned(16#24#, 8);
  gmul3_15(28) <= to_unsigned(16#27#, 8);
  gmul3_15(29) <= to_unsigned(16#22#, 8);
  gmul3_15(30) <= to_unsigned(16#21#, 8);
  gmul3_15(31) <= to_unsigned(16#60#, 8);
  gmul3_15(32) <= to_unsigned(16#63#, 8);
  gmul3_15(33) <= to_unsigned(16#66#, 8);
  gmul3_15(34) <= to_unsigned(16#65#, 8);
  gmul3_15(35) <= to_unsigned(16#6C#, 8);
  gmul3_15(36) <= to_unsigned(16#6F#, 8);
  gmul3_15(37) <= to_unsigned(16#6A#, 8);
  gmul3_15(38) <= to_unsigned(16#69#, 8);
  gmul3_15(39) <= to_unsigned(16#78#, 8);
  gmul3_15(40) <= to_unsigned(16#7B#, 8);
  gmul3_15(41) <= to_unsigned(16#7E#, 8);
  gmul3_15(42) <= to_unsigned(16#7D#, 8);
  gmul3_15(43) <= to_unsigned(16#74#, 8);
  gmul3_15(44) <= to_unsigned(16#77#, 8);
  gmul3_15(45) <= to_unsigned(16#72#, 8);
  gmul3_15(46) <= to_unsigned(16#71#, 8);
  gmul3_15(47) <= to_unsigned(16#50#, 8);
  gmul3_15(48) <= to_unsigned(16#53#, 8);
  gmul3_15(49) <= to_unsigned(16#56#, 8);
  gmul3_15(50) <= to_unsigned(16#55#, 8);
  gmul3_15(51) <= to_unsigned(16#5C#, 8);
  gmul3_15(52) <= to_unsigned(16#5F#, 8);
  gmul3_15(53) <= to_unsigned(16#5A#, 8);
  gmul3_15(54) <= to_unsigned(16#59#, 8);
  gmul3_15(55) <= to_unsigned(16#48#, 8);
  gmul3_15(56) <= to_unsigned(16#4B#, 8);
  gmul3_15(57) <= to_unsigned(16#4E#, 8);
  gmul3_15(58) <= to_unsigned(16#4D#, 8);
  gmul3_15(59) <= to_unsigned(16#44#, 8);
  gmul3_15(60) <= to_unsigned(16#47#, 8);
  gmul3_15(61) <= to_unsigned(16#42#, 8);
  gmul3_15(62) <= to_unsigned(16#41#, 8);
  gmul3_15(63) <= to_unsigned(16#C0#, 8);
  gmul3_15(64) <= to_unsigned(16#C3#, 8);
  gmul3_15(65) <= to_unsigned(16#C6#, 8);
  gmul3_15(66) <= to_unsigned(16#C5#, 8);
  gmul3_15(67) <= to_unsigned(16#CC#, 8);
  gmul3_15(68) <= to_unsigned(16#CF#, 8);
  gmul3_15(69) <= to_unsigned(16#CA#, 8);
  gmul3_15(70) <= to_unsigned(16#C9#, 8);
  gmul3_15(71) <= to_unsigned(16#D8#, 8);
  gmul3_15(72) <= to_unsigned(16#DB#, 8);
  gmul3_15(73) <= to_unsigned(16#DE#, 8);
  gmul3_15(74) <= to_unsigned(16#DD#, 8);
  gmul3_15(75) <= to_unsigned(16#D4#, 8);
  gmul3_15(76) <= to_unsigned(16#D7#, 8);
  gmul3_15(77) <= to_unsigned(16#D2#, 8);
  gmul3_15(78) <= to_unsigned(16#D1#, 8);
  gmul3_15(79) <= to_unsigned(16#F0#, 8);
  gmul3_15(80) <= to_unsigned(16#F3#, 8);
  gmul3_15(81) <= to_unsigned(16#F6#, 8);
  gmul3_15(82) <= to_unsigned(16#F5#, 8);
  gmul3_15(83) <= to_unsigned(16#FC#, 8);
  gmul3_15(84) <= to_unsigned(16#FF#, 8);
  gmul3_15(85) <= to_unsigned(16#FA#, 8);
  gmul3_15(86) <= to_unsigned(16#F9#, 8);
  gmul3_15(87) <= to_unsigned(16#E8#, 8);
  gmul3_15(88) <= to_unsigned(16#EB#, 8);
  gmul3_15(89) <= to_unsigned(16#EE#, 8);
  gmul3_15(90) <= to_unsigned(16#ED#, 8);
  gmul3_15(91) <= to_unsigned(16#E4#, 8);
  gmul3_15(92) <= to_unsigned(16#E7#, 8);
  gmul3_15(93) <= to_unsigned(16#E2#, 8);
  gmul3_15(94) <= to_unsigned(16#E1#, 8);
  gmul3_15(95) <= to_unsigned(16#A0#, 8);
  gmul3_15(96) <= to_unsigned(16#A3#, 8);
  gmul3_15(97) <= to_unsigned(16#A6#, 8);
  gmul3_15(98) <= to_unsigned(16#A5#, 8);
  gmul3_15(99) <= to_unsigned(16#AC#, 8);
  gmul3_15(100) <= to_unsigned(16#AF#, 8);
  gmul3_15(101) <= to_unsigned(16#AA#, 8);
  gmul3_15(102) <= to_unsigned(16#A9#, 8);
  gmul3_15(103) <= to_unsigned(16#B8#, 8);
  gmul3_15(104) <= to_unsigned(16#BB#, 8);
  gmul3_15(105) <= to_unsigned(16#BE#, 8);
  gmul3_15(106) <= to_unsigned(16#BD#, 8);
  gmul3_15(107) <= to_unsigned(16#B4#, 8);
  gmul3_15(108) <= to_unsigned(16#B7#, 8);
  gmul3_15(109) <= to_unsigned(16#B2#, 8);
  gmul3_15(110) <= to_unsigned(16#B1#, 8);
  gmul3_15(111) <= to_unsigned(16#90#, 8);
  gmul3_15(112) <= to_unsigned(16#93#, 8);
  gmul3_15(113) <= to_unsigned(16#96#, 8);
  gmul3_15(114) <= to_unsigned(16#95#, 8);
  gmul3_15(115) <= to_unsigned(16#9C#, 8);
  gmul3_15(116) <= to_unsigned(16#9F#, 8);
  gmul3_15(117) <= to_unsigned(16#9A#, 8);
  gmul3_15(118) <= to_unsigned(16#99#, 8);
  gmul3_15(119) <= to_unsigned(16#88#, 8);
  gmul3_15(120) <= to_unsigned(16#8B#, 8);
  gmul3_15(121) <= to_unsigned(16#8E#, 8);
  gmul3_15(122) <= to_unsigned(16#8D#, 8);
  gmul3_15(123) <= to_unsigned(16#84#, 8);
  gmul3_15(124) <= to_unsigned(16#87#, 8);
  gmul3_15(125) <= to_unsigned(16#82#, 8);
  gmul3_15(126) <= to_unsigned(16#81#, 8);
  gmul3_15(127) <= to_unsigned(16#9B#, 8);
  gmul3_15(128) <= to_unsigned(16#98#, 8);
  gmul3_15(129) <= to_unsigned(16#9D#, 8);
  gmul3_15(130) <= to_unsigned(16#9E#, 8);
  gmul3_15(131) <= to_unsigned(16#97#, 8);
  gmul3_15(132) <= to_unsigned(16#94#, 8);
  gmul3_15(133) <= to_unsigned(16#91#, 8);
  gmul3_15(134) <= to_unsigned(16#92#, 8);
  gmul3_15(135) <= to_unsigned(16#83#, 8);
  gmul3_15(136) <= to_unsigned(16#80#, 8);
  gmul3_15(137) <= to_unsigned(16#85#, 8);
  gmul3_15(138) <= to_unsigned(16#86#, 8);
  gmul3_15(139) <= to_unsigned(16#8F#, 8);
  gmul3_15(140) <= to_unsigned(16#8C#, 8);
  gmul3_15(141) <= to_unsigned(16#89#, 8);
  gmul3_15(142) <= to_unsigned(16#8A#, 8);
  gmul3_15(143) <= to_unsigned(16#AB#, 8);
  gmul3_15(144) <= to_unsigned(16#A8#, 8);
  gmul3_15(145) <= to_unsigned(16#AD#, 8);
  gmul3_15(146) <= to_unsigned(16#AE#, 8);
  gmul3_15(147) <= to_unsigned(16#A7#, 8);
  gmul3_15(148) <= to_unsigned(16#A4#, 8);
  gmul3_15(149) <= to_unsigned(16#A1#, 8);
  gmul3_15(150) <= to_unsigned(16#A2#, 8);
  gmul3_15(151) <= to_unsigned(16#B3#, 8);
  gmul3_15(152) <= to_unsigned(16#B0#, 8);
  gmul3_15(153) <= to_unsigned(16#B5#, 8);
  gmul3_15(154) <= to_unsigned(16#B6#, 8);
  gmul3_15(155) <= to_unsigned(16#BF#, 8);
  gmul3_15(156) <= to_unsigned(16#BC#, 8);
  gmul3_15(157) <= to_unsigned(16#B9#, 8);
  gmul3_15(158) <= to_unsigned(16#BA#, 8);
  gmul3_15(159) <= to_unsigned(16#FB#, 8);
  gmul3_15(160) <= to_unsigned(16#F8#, 8);
  gmul3_15(161) <= to_unsigned(16#FD#, 8);
  gmul3_15(162) <= to_unsigned(16#FE#, 8);
  gmul3_15(163) <= to_unsigned(16#F7#, 8);
  gmul3_15(164) <= to_unsigned(16#F4#, 8);
  gmul3_15(165) <= to_unsigned(16#F1#, 8);
  gmul3_15(166) <= to_unsigned(16#F2#, 8);
  gmul3_15(167) <= to_unsigned(16#E3#, 8);
  gmul3_15(168) <= to_unsigned(16#E0#, 8);
  gmul3_15(169) <= to_unsigned(16#E5#, 8);
  gmul3_15(170) <= to_unsigned(16#E6#, 8);
  gmul3_15(171) <= to_unsigned(16#EF#, 8);
  gmul3_15(172) <= to_unsigned(16#EC#, 8);
  gmul3_15(173) <= to_unsigned(16#E9#, 8);
  gmul3_15(174) <= to_unsigned(16#EA#, 8);
  gmul3_15(175) <= to_unsigned(16#CB#, 8);
  gmul3_15(176) <= to_unsigned(16#C8#, 8);
  gmul3_15(177) <= to_unsigned(16#CD#, 8);
  gmul3_15(178) <= to_unsigned(16#CE#, 8);
  gmul3_15(179) <= to_unsigned(16#C7#, 8);
  gmul3_15(180) <= to_unsigned(16#C4#, 8);
  gmul3_15(181) <= to_unsigned(16#C1#, 8);
  gmul3_15(182) <= to_unsigned(16#C2#, 8);
  gmul3_15(183) <= to_unsigned(16#D3#, 8);
  gmul3_15(184) <= to_unsigned(16#D0#, 8);
  gmul3_15(185) <= to_unsigned(16#D5#, 8);
  gmul3_15(186) <= to_unsigned(16#D6#, 8);
  gmul3_15(187) <= to_unsigned(16#DF#, 8);
  gmul3_15(188) <= to_unsigned(16#DC#, 8);
  gmul3_15(189) <= to_unsigned(16#D9#, 8);
  gmul3_15(190) <= to_unsigned(16#DA#, 8);
  gmul3_15(191) <= to_unsigned(16#5B#, 8);
  gmul3_15(192) <= to_unsigned(16#58#, 8);
  gmul3_15(193) <= to_unsigned(16#5D#, 8);
  gmul3_15(194) <= to_unsigned(16#5E#, 8);
  gmul3_15(195) <= to_unsigned(16#57#, 8);
  gmul3_15(196) <= to_unsigned(16#54#, 8);
  gmul3_15(197) <= to_unsigned(16#51#, 8);
  gmul3_15(198) <= to_unsigned(16#52#, 8);
  gmul3_15(199) <= to_unsigned(16#43#, 8);
  gmul3_15(200) <= to_unsigned(16#40#, 8);
  gmul3_15(201) <= to_unsigned(16#45#, 8);
  gmul3_15(202) <= to_unsigned(16#46#, 8);
  gmul3_15(203) <= to_unsigned(16#4F#, 8);
  gmul3_15(204) <= to_unsigned(16#4C#, 8);
  gmul3_15(205) <= to_unsigned(16#49#, 8);
  gmul3_15(206) <= to_unsigned(16#4A#, 8);
  gmul3_15(207) <= to_unsigned(16#6B#, 8);
  gmul3_15(208) <= to_unsigned(16#68#, 8);
  gmul3_15(209) <= to_unsigned(16#6D#, 8);
  gmul3_15(210) <= to_unsigned(16#6E#, 8);
  gmul3_15(211) <= to_unsigned(16#67#, 8);
  gmul3_15(212) <= to_unsigned(16#64#, 8);
  gmul3_15(213) <= to_unsigned(16#61#, 8);
  gmul3_15(214) <= to_unsigned(16#62#, 8);
  gmul3_15(215) <= to_unsigned(16#73#, 8);
  gmul3_15(216) <= to_unsigned(16#70#, 8);
  gmul3_15(217) <= to_unsigned(16#75#, 8);
  gmul3_15(218) <= to_unsigned(16#76#, 8);
  gmul3_15(219) <= to_unsigned(16#7F#, 8);
  gmul3_15(220) <= to_unsigned(16#7C#, 8);
  gmul3_15(221) <= to_unsigned(16#79#, 8);
  gmul3_15(222) <= to_unsigned(16#7A#, 8);
  gmul3_15(223) <= to_unsigned(16#3B#, 8);
  gmul3_15(224) <= to_unsigned(16#38#, 8);
  gmul3_15(225) <= to_unsigned(16#3D#, 8);
  gmul3_15(226) <= to_unsigned(16#3E#, 8);
  gmul3_15(227) <= to_unsigned(16#37#, 8);
  gmul3_15(228) <= to_unsigned(16#34#, 8);
  gmul3_15(229) <= to_unsigned(16#31#, 8);
  gmul3_15(230) <= to_unsigned(16#32#, 8);
  gmul3_15(231) <= to_unsigned(16#23#, 8);
  gmul3_15(232) <= to_unsigned(16#20#, 8);
  gmul3_15(233) <= to_unsigned(16#25#, 8);
  gmul3_15(234) <= to_unsigned(16#26#, 8);
  gmul3_15(235) <= to_unsigned(16#2F#, 8);
  gmul3_15(236) <= to_unsigned(16#2C#, 8);
  gmul3_15(237) <= to_unsigned(16#29#, 8);
  gmul3_15(238) <= to_unsigned(16#2A#, 8);
  gmul3_15(239) <= to_unsigned(16#0B#, 8);
  gmul3_15(240) <= to_unsigned(16#08#, 8);
  gmul3_15(241) <= to_unsigned(16#0D#, 8);
  gmul3_15(242) <= to_unsigned(16#0E#, 8);
  gmul3_15(243) <= to_unsigned(16#07#, 8);
  gmul3_15(244) <= to_unsigned(16#04#, 8);
  gmul3_15(245) <= to_unsigned(16#01#, 8);
  gmul3_15(246) <= to_unsigned(16#02#, 8);
  gmul3_15(247) <= to_unsigned(16#13#, 8);
  gmul3_15(248) <= to_unsigned(16#10#, 8);
  gmul3_15(249) <= to_unsigned(16#15#, 8);
  gmul3_15(250) <= to_unsigned(16#16#, 8);
  gmul3_15(251) <= to_unsigned(16#1F#, 8);
  gmul3_15(252) <= to_unsigned(16#1C#, 8);
  gmul3_15(253) <= to_unsigned(16#19#, 8);
  gmul3_15(254) <= to_unsigned(16#1A#, 8);
  gmul3_15(255) <= to_unsigned(16#1A#, 8);

  gmul2_15(0) <= to_unsigned(16#02#, 8);
  gmul2_15(1) <= to_unsigned(16#04#, 8);
  gmul2_15(2) <= to_unsigned(16#06#, 8);
  gmul2_15(3) <= to_unsigned(16#08#, 8);
  gmul2_15(4) <= to_unsigned(16#0A#, 8);
  gmul2_15(5) <= to_unsigned(16#0C#, 8);
  gmul2_15(6) <= to_unsigned(16#0E#, 8);
  gmul2_15(7) <= to_unsigned(16#10#, 8);
  gmul2_15(8) <= to_unsigned(16#12#, 8);
  gmul2_15(9) <= to_unsigned(16#14#, 8);
  gmul2_15(10) <= to_unsigned(16#16#, 8);
  gmul2_15(11) <= to_unsigned(16#18#, 8);
  gmul2_15(12) <= to_unsigned(16#1A#, 8);
  gmul2_15(13) <= to_unsigned(16#1C#, 8);
  gmul2_15(14) <= to_unsigned(16#1E#, 8);
  gmul2_15(15) <= to_unsigned(16#20#, 8);
  gmul2_15(16) <= to_unsigned(16#22#, 8);
  gmul2_15(17) <= to_unsigned(16#24#, 8);
  gmul2_15(18) <= to_unsigned(16#26#, 8);
  gmul2_15(19) <= to_unsigned(16#28#, 8);
  gmul2_15(20) <= to_unsigned(16#2A#, 8);
  gmul2_15(21) <= to_unsigned(16#2C#, 8);
  gmul2_15(22) <= to_unsigned(16#2E#, 8);
  gmul2_15(23) <= to_unsigned(16#30#, 8);
  gmul2_15(24) <= to_unsigned(16#32#, 8);
  gmul2_15(25) <= to_unsigned(16#34#, 8);
  gmul2_15(26) <= to_unsigned(16#36#, 8);
  gmul2_15(27) <= to_unsigned(16#38#, 8);
  gmul2_15(28) <= to_unsigned(16#3A#, 8);
  gmul2_15(29) <= to_unsigned(16#3C#, 8);
  gmul2_15(30) <= to_unsigned(16#3E#, 8);
  gmul2_15(31) <= to_unsigned(16#40#, 8);
  gmul2_15(32) <= to_unsigned(16#42#, 8);
  gmul2_15(33) <= to_unsigned(16#44#, 8);
  gmul2_15(34) <= to_unsigned(16#46#, 8);
  gmul2_15(35) <= to_unsigned(16#48#, 8);
  gmul2_15(36) <= to_unsigned(16#4A#, 8);
  gmul2_15(37) <= to_unsigned(16#4C#, 8);
  gmul2_15(38) <= to_unsigned(16#4E#, 8);
  gmul2_15(39) <= to_unsigned(16#50#, 8);
  gmul2_15(40) <= to_unsigned(16#52#, 8);
  gmul2_15(41) <= to_unsigned(16#54#, 8);
  gmul2_15(42) <= to_unsigned(16#56#, 8);
  gmul2_15(43) <= to_unsigned(16#58#, 8);
  gmul2_15(44) <= to_unsigned(16#5A#, 8);
  gmul2_15(45) <= to_unsigned(16#5C#, 8);
  gmul2_15(46) <= to_unsigned(16#5E#, 8);
  gmul2_15(47) <= to_unsigned(16#60#, 8);
  gmul2_15(48) <= to_unsigned(16#62#, 8);
  gmul2_15(49) <= to_unsigned(16#64#, 8);
  gmul2_15(50) <= to_unsigned(16#66#, 8);
  gmul2_15(51) <= to_unsigned(16#68#, 8);
  gmul2_15(52) <= to_unsigned(16#6A#, 8);
  gmul2_15(53) <= to_unsigned(16#6C#, 8);
  gmul2_15(54) <= to_unsigned(16#6E#, 8);
  gmul2_15(55) <= to_unsigned(16#70#, 8);
  gmul2_15(56) <= to_unsigned(16#72#, 8);
  gmul2_15(57) <= to_unsigned(16#74#, 8);
  gmul2_15(58) <= to_unsigned(16#76#, 8);
  gmul2_15(59) <= to_unsigned(16#78#, 8);
  gmul2_15(60) <= to_unsigned(16#7A#, 8);
  gmul2_15(61) <= to_unsigned(16#7C#, 8);
  gmul2_15(62) <= to_unsigned(16#7E#, 8);
  gmul2_15(63) <= to_unsigned(16#80#, 8);
  gmul2_15(64) <= to_unsigned(16#82#, 8);
  gmul2_15(65) <= to_unsigned(16#84#, 8);
  gmul2_15(66) <= to_unsigned(16#86#, 8);
  gmul2_15(67) <= to_unsigned(16#88#, 8);
  gmul2_15(68) <= to_unsigned(16#8A#, 8);
  gmul2_15(69) <= to_unsigned(16#8C#, 8);
  gmul2_15(70) <= to_unsigned(16#8E#, 8);
  gmul2_15(71) <= to_unsigned(16#90#, 8);
  gmul2_15(72) <= to_unsigned(16#92#, 8);
  gmul2_15(73) <= to_unsigned(16#94#, 8);
  gmul2_15(74) <= to_unsigned(16#96#, 8);
  gmul2_15(75) <= to_unsigned(16#98#, 8);
  gmul2_15(76) <= to_unsigned(16#9A#, 8);
  gmul2_15(77) <= to_unsigned(16#9C#, 8);
  gmul2_15(78) <= to_unsigned(16#9E#, 8);
  gmul2_15(79) <= to_unsigned(16#A0#, 8);
  gmul2_15(80) <= to_unsigned(16#A2#, 8);
  gmul2_15(81) <= to_unsigned(16#A4#, 8);
  gmul2_15(82) <= to_unsigned(16#A6#, 8);
  gmul2_15(83) <= to_unsigned(16#A8#, 8);
  gmul2_15(84) <= to_unsigned(16#AA#, 8);
  gmul2_15(85) <= to_unsigned(16#AC#, 8);
  gmul2_15(86) <= to_unsigned(16#AE#, 8);
  gmul2_15(87) <= to_unsigned(16#B0#, 8);
  gmul2_15(88) <= to_unsigned(16#B2#, 8);
  gmul2_15(89) <= to_unsigned(16#B4#, 8);
  gmul2_15(90) <= to_unsigned(16#B6#, 8);
  gmul2_15(91) <= to_unsigned(16#B8#, 8);
  gmul2_15(92) <= to_unsigned(16#BA#, 8);
  gmul2_15(93) <= to_unsigned(16#BC#, 8);
  gmul2_15(94) <= to_unsigned(16#BE#, 8);
  gmul2_15(95) <= to_unsigned(16#C0#, 8);
  gmul2_15(96) <= to_unsigned(16#C2#, 8);
  gmul2_15(97) <= to_unsigned(16#C4#, 8);
  gmul2_15(98) <= to_unsigned(16#C6#, 8);
  gmul2_15(99) <= to_unsigned(16#C8#, 8);
  gmul2_15(100) <= to_unsigned(16#CA#, 8);
  gmul2_15(101) <= to_unsigned(16#CC#, 8);
  gmul2_15(102) <= to_unsigned(16#CE#, 8);
  gmul2_15(103) <= to_unsigned(16#D0#, 8);
  gmul2_15(104) <= to_unsigned(16#D2#, 8);
  gmul2_15(105) <= to_unsigned(16#D4#, 8);
  gmul2_15(106) <= to_unsigned(16#D6#, 8);
  gmul2_15(107) <= to_unsigned(16#D8#, 8);
  gmul2_15(108) <= to_unsigned(16#DA#, 8);
  gmul2_15(109) <= to_unsigned(16#DC#, 8);
  gmul2_15(110) <= to_unsigned(16#DE#, 8);
  gmul2_15(111) <= to_unsigned(16#E0#, 8);
  gmul2_15(112) <= to_unsigned(16#E2#, 8);
  gmul2_15(113) <= to_unsigned(16#E4#, 8);
  gmul2_15(114) <= to_unsigned(16#E6#, 8);
  gmul2_15(115) <= to_unsigned(16#E8#, 8);
  gmul2_15(116) <= to_unsigned(16#EA#, 8);
  gmul2_15(117) <= to_unsigned(16#EC#, 8);
  gmul2_15(118) <= to_unsigned(16#EE#, 8);
  gmul2_15(119) <= to_unsigned(16#F0#, 8);
  gmul2_15(120) <= to_unsigned(16#F2#, 8);
  gmul2_15(121) <= to_unsigned(16#F4#, 8);
  gmul2_15(122) <= to_unsigned(16#F6#, 8);
  gmul2_15(123) <= to_unsigned(16#F8#, 8);
  gmul2_15(124) <= to_unsigned(16#FA#, 8);
  gmul2_15(125) <= to_unsigned(16#FC#, 8);
  gmul2_15(126) <= to_unsigned(16#FE#, 8);
  gmul2_15(127) <= to_unsigned(16#1B#, 8);
  gmul2_15(128) <= to_unsigned(16#19#, 8);
  gmul2_15(129) <= to_unsigned(16#1F#, 8);
  gmul2_15(130) <= to_unsigned(16#1D#, 8);
  gmul2_15(131) <= to_unsigned(16#13#, 8);
  gmul2_15(132) <= to_unsigned(16#11#, 8);
  gmul2_15(133) <= to_unsigned(16#17#, 8);
  gmul2_15(134) <= to_unsigned(16#15#, 8);
  gmul2_15(135) <= to_unsigned(16#0B#, 8);
  gmul2_15(136) <= to_unsigned(16#09#, 8);
  gmul2_15(137) <= to_unsigned(16#0F#, 8);
  gmul2_15(138) <= to_unsigned(16#0D#, 8);
  gmul2_15(139) <= to_unsigned(16#03#, 8);
  gmul2_15(140) <= to_unsigned(16#01#, 8);
  gmul2_15(141) <= to_unsigned(16#07#, 8);
  gmul2_15(142) <= to_unsigned(16#05#, 8);
  gmul2_15(143) <= to_unsigned(16#3B#, 8);
  gmul2_15(144) <= to_unsigned(16#39#, 8);
  gmul2_15(145) <= to_unsigned(16#3F#, 8);
  gmul2_15(146) <= to_unsigned(16#3D#, 8);
  gmul2_15(147) <= to_unsigned(16#33#, 8);
  gmul2_15(148) <= to_unsigned(16#31#, 8);
  gmul2_15(149) <= to_unsigned(16#37#, 8);
  gmul2_15(150) <= to_unsigned(16#35#, 8);
  gmul2_15(151) <= to_unsigned(16#2B#, 8);
  gmul2_15(152) <= to_unsigned(16#29#, 8);
  gmul2_15(153) <= to_unsigned(16#2F#, 8);
  gmul2_15(154) <= to_unsigned(16#2D#, 8);
  gmul2_15(155) <= to_unsigned(16#23#, 8);
  gmul2_15(156) <= to_unsigned(16#21#, 8);
  gmul2_15(157) <= to_unsigned(16#27#, 8);
  gmul2_15(158) <= to_unsigned(16#25#, 8);
  gmul2_15(159) <= to_unsigned(16#5B#, 8);
  gmul2_15(160) <= to_unsigned(16#59#, 8);
  gmul2_15(161) <= to_unsigned(16#5F#, 8);
  gmul2_15(162) <= to_unsigned(16#5D#, 8);
  gmul2_15(163) <= to_unsigned(16#53#, 8);
  gmul2_15(164) <= to_unsigned(16#51#, 8);
  gmul2_15(165) <= to_unsigned(16#57#, 8);
  gmul2_15(166) <= to_unsigned(16#55#, 8);
  gmul2_15(167) <= to_unsigned(16#4B#, 8);
  gmul2_15(168) <= to_unsigned(16#49#, 8);
  gmul2_15(169) <= to_unsigned(16#4F#, 8);
  gmul2_15(170) <= to_unsigned(16#4D#, 8);
  gmul2_15(171) <= to_unsigned(16#43#, 8);
  gmul2_15(172) <= to_unsigned(16#41#, 8);
  gmul2_15(173) <= to_unsigned(16#47#, 8);
  gmul2_15(174) <= to_unsigned(16#45#, 8);
  gmul2_15(175) <= to_unsigned(16#7B#, 8);
  gmul2_15(176) <= to_unsigned(16#79#, 8);
  gmul2_15(177) <= to_unsigned(16#7F#, 8);
  gmul2_15(178) <= to_unsigned(16#7D#, 8);
  gmul2_15(179) <= to_unsigned(16#73#, 8);
  gmul2_15(180) <= to_unsigned(16#71#, 8);
  gmul2_15(181) <= to_unsigned(16#77#, 8);
  gmul2_15(182) <= to_unsigned(16#75#, 8);
  gmul2_15(183) <= to_unsigned(16#6B#, 8);
  gmul2_15(184) <= to_unsigned(16#69#, 8);
  gmul2_15(185) <= to_unsigned(16#6F#, 8);
  gmul2_15(186) <= to_unsigned(16#6D#, 8);
  gmul2_15(187) <= to_unsigned(16#63#, 8);
  gmul2_15(188) <= to_unsigned(16#61#, 8);
  gmul2_15(189) <= to_unsigned(16#67#, 8);
  gmul2_15(190) <= to_unsigned(16#65#, 8);
  gmul2_15(191) <= to_unsigned(16#9B#, 8);
  gmul2_15(192) <= to_unsigned(16#99#, 8);
  gmul2_15(193) <= to_unsigned(16#9F#, 8);
  gmul2_15(194) <= to_unsigned(16#9D#, 8);
  gmul2_15(195) <= to_unsigned(16#93#, 8);
  gmul2_15(196) <= to_unsigned(16#91#, 8);
  gmul2_15(197) <= to_unsigned(16#97#, 8);
  gmul2_15(198) <= to_unsigned(16#95#, 8);
  gmul2_15(199) <= to_unsigned(16#8B#, 8);
  gmul2_15(200) <= to_unsigned(16#89#, 8);
  gmul2_15(201) <= to_unsigned(16#8F#, 8);
  gmul2_15(202) <= to_unsigned(16#8D#, 8);
  gmul2_15(203) <= to_unsigned(16#83#, 8);
  gmul2_15(204) <= to_unsigned(16#81#, 8);
  gmul2_15(205) <= to_unsigned(16#87#, 8);
  gmul2_15(206) <= to_unsigned(16#85#, 8);
  gmul2_15(207) <= to_unsigned(16#BB#, 8);
  gmul2_15(208) <= to_unsigned(16#B9#, 8);
  gmul2_15(209) <= to_unsigned(16#BF#, 8);
  gmul2_15(210) <= to_unsigned(16#BD#, 8);
  gmul2_15(211) <= to_unsigned(16#B3#, 8);
  gmul2_15(212) <= to_unsigned(16#B1#, 8);
  gmul2_15(213) <= to_unsigned(16#B7#, 8);
  gmul2_15(214) <= to_unsigned(16#B5#, 8);
  gmul2_15(215) <= to_unsigned(16#AB#, 8);
  gmul2_15(216) <= to_unsigned(16#A9#, 8);
  gmul2_15(217) <= to_unsigned(16#AF#, 8);
  gmul2_15(218) <= to_unsigned(16#AD#, 8);
  gmul2_15(219) <= to_unsigned(16#A3#, 8);
  gmul2_15(220) <= to_unsigned(16#A1#, 8);
  gmul2_15(221) <= to_unsigned(16#A7#, 8);
  gmul2_15(222) <= to_unsigned(16#A5#, 8);
  gmul2_15(223) <= to_unsigned(16#DB#, 8);
  gmul2_15(224) <= to_unsigned(16#D9#, 8);
  gmul2_15(225) <= to_unsigned(16#DF#, 8);
  gmul2_15(226) <= to_unsigned(16#DD#, 8);
  gmul2_15(227) <= to_unsigned(16#D3#, 8);
  gmul2_15(228) <= to_unsigned(16#D1#, 8);
  gmul2_15(229) <= to_unsigned(16#D7#, 8);
  gmul2_15(230) <= to_unsigned(16#D5#, 8);
  gmul2_15(231) <= to_unsigned(16#CB#, 8);
  gmul2_15(232) <= to_unsigned(16#C9#, 8);
  gmul2_15(233) <= to_unsigned(16#CF#, 8);
  gmul2_15(234) <= to_unsigned(16#CD#, 8);
  gmul2_15(235) <= to_unsigned(16#C3#, 8);
  gmul2_15(236) <= to_unsigned(16#C1#, 8);
  gmul2_15(237) <= to_unsigned(16#C7#, 8);
  gmul2_15(238) <= to_unsigned(16#C5#, 8);
  gmul2_15(239) <= to_unsigned(16#FB#, 8);
  gmul2_15(240) <= to_unsigned(16#F9#, 8);
  gmul2_15(241) <= to_unsigned(16#FF#, 8);
  gmul2_15(242) <= to_unsigned(16#FD#, 8);
  gmul2_15(243) <= to_unsigned(16#F3#, 8);
  gmul2_15(244) <= to_unsigned(16#F1#, 8);
  gmul2_15(245) <= to_unsigned(16#F7#, 8);
  gmul2_15(246) <= to_unsigned(16#F5#, 8);
  gmul2_15(247) <= to_unsigned(16#EB#, 8);
  gmul2_15(248) <= to_unsigned(16#E9#, 8);
  gmul2_15(249) <= to_unsigned(16#EF#, 8);
  gmul2_15(250) <= to_unsigned(16#ED#, 8);
  gmul2_15(251) <= to_unsigned(16#E3#, 8);
  gmul2_15(252) <= to_unsigned(16#E1#, 8);
  gmul2_15(253) <= to_unsigned(16#E7#, 8);
  gmul2_15(254) <= to_unsigned(16#E5#, 8);
  gmul2_15(255) <= to_unsigned(16#E5#, 8);

  const_expression_26 <= to_unsigned(16#0001#, 16);

  out0_122(0) <= expandedKey(0);
  out0_122(1) <= expandedKey(1);
  out0_122(2) <= expandedKey(2);
  out0_122(3) <= expandedKey(3);
  out0_122(4) <= expandedKey(4);
  out0_122(5) <= expandedKey(5);
  out0_122(6) <= expandedKey(6);
  out0_122(7) <= expandedKey(7);
  out0_122(8) <= expandedKey(8);
  out0_122(9) <= expandedKey(9);
  out0_122(10) <= expandedKey(10);
  out0_122(11) <= expandedKey(11);
  out0_122(12) <= expandedKey(12);
  out0_122(13) <= expandedKey(13);
  out0_122(14) <= expandedKey(14);
  out0_122(15) <= expandedKey(15);

  inBytes_signal1_unsigned <= unsigned(inBytes_signal1);

  Delay1_1_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal1_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal1_1 <= inBytes_signal1_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_1_process;


  inBytes_signal2_unsigned <= unsigned(inBytes_signal2);

  Delay1_2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal2_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal2_1 <= inBytes_signal2_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_2_process;


  inBytes_signal3_unsigned <= unsigned(inBytes_signal3);

  Delay1_3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal3_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal3_1 <= inBytes_signal3_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_3_process;


  inBytes_signal4_unsigned <= unsigned(inBytes_signal4);

  Delay1_4_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal4_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal4_1 <= inBytes_signal4_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_4_process;


  inBytes_signal5_unsigned <= unsigned(inBytes_signal5);

  Delay1_5_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal5_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal5_1 <= inBytes_signal5_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_5_process;


  inBytes_signal6_unsigned <= unsigned(inBytes_signal6);

  Delay1_6_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal6_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal6_1 <= inBytes_signal6_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_6_process;


  inBytes_signal7_unsigned <= unsigned(inBytes_signal7);

  Delay1_7_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal7_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal7_1 <= inBytes_signal7_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_7_process;


  inBytes_signal8_unsigned <= unsigned(inBytes_signal8);

  Delay1_8_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal8_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal8_1 <= inBytes_signal8_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_8_process;


  inBytes_signal9_unsigned <= unsigned(inBytes_signal9);

  Delay1_9_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal9_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal9_1 <= inBytes_signal9_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_9_process;


  inBytes_signal10_unsigned <= unsigned(inBytes_signal10);

  Delay1_10_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal10_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal10_1 <= inBytes_signal10_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_10_process;


  inBytes_signal11_unsigned <= unsigned(inBytes_signal11);

  Delay1_11_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal11_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal11_1 <= inBytes_signal11_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_11_process;


  inBytes_signal12_unsigned <= unsigned(inBytes_signal12);

  Delay1_12_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal12_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal12_1 <= inBytes_signal12_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_12_process;


  inBytes_signal13_unsigned <= unsigned(inBytes_signal13);

  Delay1_13_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal13_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal13_1 <= inBytes_signal13_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_13_process;


  inBytes_signal14_unsigned <= unsigned(inBytes_signal14);

  Delay1_14_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal14_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal14_1 <= inBytes_signal14_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_14_process;


  inBytes_signal15_unsigned <= unsigned(inBytes_signal15);

  Delay1_15_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal15_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal15_1 <= inBytes_signal15_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_15_process;


  inBytes_signal16_unsigned <= unsigned(inBytes_signal16);

  Delay1_16_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        signal16_1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        signal16_1 <= inBytes_signal16_unsigned;
      END IF;
    END IF;
  END PROCESS Delay1_16_process;


  Delay1_out1_to_vector(0) <= signal1_1;
  Delay1_out1_to_vector(1) <= signal2_1;
  Delay1_out1_to_vector(2) <= signal3_1;
  Delay1_out1_to_vector(3) <= signal4_1;
  Delay1_out1_to_vector(4) <= signal5_1;
  Delay1_out1_to_vector(5) <= signal6_1;
  Delay1_out1_to_vector(6) <= signal7_1;
  Delay1_out1_to_vector(7) <= signal8_1;
  Delay1_out1_to_vector(8) <= signal9_1;
  Delay1_out1_to_vector(9) <= signal10_1;
  Delay1_out1_to_vector(10) <= signal11_1;
  Delay1_out1_to_vector(11) <= signal12_1;
  Delay1_out1_to_vector(12) <= signal13_1;
  Delay1_out1_to_vector(13) <= signal14_1;
  Delay1_out1_to_vector(14) <= signal15_1;
  Delay1_out1_to_vector(15) <= signal16_1;

  s_s(0) <= Delay1_out1_to_vector(0);
  s_s(1) <= Delay1_out1_to_vector(1);
  s_s(2) <= Delay1_out1_to_vector(2);
  s_s(3) <= Delay1_out1_to_vector(3);
  s_s(4) <= Delay1_out1_to_vector(4);
  s_s(5) <= Delay1_out1_to_vector(5);
  s_s(6) <= Delay1_out1_to_vector(6);
  s_s(7) <= Delay1_out1_to_vector(7);
  s_s(8) <= Delay1_out1_to_vector(8);
  s_s(9) <= Delay1_out1_to_vector(9);
  s_s(10) <= Delay1_out1_to_vector(10);
  s_s(11) <= Delay1_out1_to_vector(11);
  s_s(12) <= Delay1_out1_to_vector(12);
  s_s(13) <= Delay1_out1_to_vector(13);
  s_s(14) <= Delay1_out1_to_vector(14);
  s_s(15) <= Delay1_out1_to_vector(15);

  out0_123(0) <= s_s_1(0);
  out0_123(1) <= s_s_1(1);
  out0_123(2) <= s_s_1(2);
  out0_123(3) <= s_s_1(3);
  out0_123(4) <= s_s_1(4);
  out0_123(5) <= s_s_1(5);
  out0_123(6) <= s_s_1(6);
  out0_123(7) <= s_s_1(7);
  out0_123(8) <= s_s_1(8);
  out0_123(9) <= s_s_1(9);
  out0_123(10) <= s_s_1(10);
  out0_123(11) <= s_s_1(11);
  out0_123(12) <= s_s_1(12);
  out0_123(13) <= s_s_1(13);
  out0_123(14) <= s_s_1(14);
  out0_123(15) <= s_s_1(15);

  s_s_2(0) <= out0_123(0) XOR out0_122(0);
  s_s_2(1) <= out0_123(1) XOR out0_122(1);
  s_s_2(2) <= out0_123(2) XOR out0_122(2);
  s_s_2(3) <= out0_123(3) XOR out0_122(3);
  s_s_2(4) <= out0_123(4) XOR out0_122(4);
  s_s_2(5) <= out0_123(5) XOR out0_122(5);
  s_s_2(6) <= out0_123(6) XOR out0_122(6);
  s_s_2(7) <= out0_123(7) XOR out0_122(7);
  s_s_2(8) <= out0_123(8) XOR out0_122(8);
  s_s_2(9) <= out0_123(9) XOR out0_122(9);
  s_s_2(10) <= out0_123(10) XOR out0_122(10);
  s_s_2(11) <= out0_123(11) XOR out0_122(11);
  s_s_2(12) <= out0_123(12) XOR out0_122(12);
  s_s_2(13) <= out0_123(13) XOR out0_122(13);
  s_s_2(14) <= out0_123(14) XOR out0_122(14);
  s_s_2(15) <= out0_123(15) XOR out0_122(15);

  out0_11_1 <= out0_124(11);

  
  s_11 <= sbox(0) WHEN out0_11_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_11_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_11_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_11_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_11_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_11_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_11_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_11_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_11_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_11_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_11_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_11_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_11_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_11_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_11_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_11_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_11_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_11_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_11_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_11_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_11_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_11_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_11_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_11_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_11_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_11_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_11_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_11_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_11_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_11_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_11_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_11_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_11_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_11_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_11_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_11_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_11_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_11_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_11_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_11_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_11_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_11_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_11_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_11_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_11_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_11_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_11_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_11_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_11_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_11_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_11_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_11_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_11_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_11_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_11_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_11_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_11_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_11_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_11_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_11_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_11_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_11_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_11_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_11_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_11_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_11_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_11_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_11_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_11_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_11_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_11_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_11_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_11_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_11_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_11_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_11_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_11_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_11_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_11_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_11_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_11_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_11_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_11_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_11_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_11_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_11_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_11_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_11_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_11_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_11_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_11_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_11_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_11_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_11_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_11_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_11_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_11_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_11_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_11_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_11_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_11_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_11_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_11_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_11_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_11_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_11_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_11_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_11_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_11_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_11_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_11_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_11_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_11_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_11_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_11_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_11_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_11_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_11_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_11_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_11_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_11_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_11_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_11_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_11_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_11_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_11_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_11_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_11_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_11_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_11_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_11_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_11_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_11_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_11_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_11_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_11_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_11_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_11_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_11_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_11_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_11_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_11_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_11_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_11_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_11_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_11_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_11_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_11_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_11_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_11_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_11_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_11_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_11_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_11_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_11_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_11_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_11_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_11_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_11_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_11_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_11_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_11_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_11_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_11_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_11_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_11_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_11_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_11_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_11_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_11_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_11_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_11_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_11_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_11_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_11_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_11_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_11_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_11_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_11_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_11_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_11_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_11_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_11_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_11_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_11_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_11_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_11_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_11_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_11_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_11_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_11_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_11_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_11_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_11_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_11_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_11_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_11_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_11_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_11_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_11_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_11_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_11_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_11_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_11_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_11_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_11_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_11_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_11_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_11_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_11_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_11_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_11_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_11_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_11_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_11_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_11_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_11_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_11_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_11_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_11_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_11_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_11_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_11_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_11_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_11_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_11_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_11_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_11_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_11_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_11_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_11_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_11_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_11_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_11_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_11_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_11_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_11_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_11_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_11_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_11_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_11_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_11_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_11_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_11_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_11_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_11_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_11_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_11_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_11_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_11_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_11_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_11_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_11_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_11_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_11_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_6_1 <= out0_124(6);

  
  s_6 <= sbox(0) WHEN out0_6_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_6_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_6_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_6_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_6_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_6_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_6_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_6_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_6_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_6_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_6_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_6_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_6_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_6_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_6_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_6_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_6_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_6_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_6_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_6_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_6_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_6_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_6_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_6_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_6_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_6_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_6_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_6_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_6_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_6_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_6_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_6_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_6_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_6_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_6_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_6_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_6_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_6_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_6_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_6_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_6_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_6_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_6_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_6_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_6_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_6_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_6_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_6_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_6_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_6_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_6_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_6_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_6_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_6_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_6_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_6_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_6_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_6_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_6_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_6_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_6_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_6_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_6_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_6_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_6_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_6_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_6_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_6_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_6_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_6_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_6_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_6_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_6_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_6_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_6_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_6_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_6_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_6_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_6_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_6_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_6_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_6_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_6_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_6_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_6_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_6_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_6_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_6_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_6_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_6_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_6_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_6_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_6_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_6_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_6_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_6_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_6_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_6_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_6_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_6_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_6_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_6_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_6_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_6_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_6_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_6_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_6_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_6_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_6_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_6_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_6_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_6_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_6_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_6_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_6_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_6_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_6_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_6_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_6_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_6_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_6_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_6_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_6_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_6_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_6_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_6_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_6_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_6_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_6_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_6_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_6_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_6_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_6_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_6_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_6_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_6_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_6_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_6_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_6_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_6_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_6_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_6_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_6_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_6_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_6_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_6_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_6_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_6_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_6_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_6_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_6_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_6_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_6_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_6_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_6_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_6_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_6_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_6_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_6_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_6_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_6_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_6_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_6_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_6_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_6_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_6_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_6_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_6_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_6_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_6_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_6_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_6_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_6_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_6_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_6_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_6_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_6_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_6_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_6_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_6_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_6_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_6_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_6_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_6_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_6_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_6_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_6_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_6_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_6_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_6_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_6_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_6_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_6_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_6_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_6_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_6_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_6_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_6_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_6_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_6_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_6_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_6_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_6_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_6_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_6_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_6_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_6_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_6_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_6_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_6_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_6_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_6_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_6_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_6_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_6_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_6_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_6_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_6_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_6_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_6_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_6_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_6_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_6_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_6_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_6_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_6_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_6_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_6_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_6_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_6_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_6_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_6_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_6_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_6_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_6_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_6_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_6_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_6_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_6_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_6_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_6_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_6_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_6_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_6_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_6_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_6_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_6_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_6_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_6_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_6_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_6_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_6_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_6_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_6_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_6_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_1_3 <= out0_124(1);

  
  s_1 <= sbox(0) WHEN out0_1_3 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_1_3 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_1_3 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_1_3 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_1_3 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_1_3 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_1_3 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_1_3 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_1_3 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_1_3 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_1_3 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_1_3 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_1_3 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_1_3 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_1_3 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_1_3 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_1_3 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_1_3 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_1_3 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_1_3 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_1_3 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_1_3 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_1_3 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_1_3 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_1_3 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_1_3 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_1_3 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_1_3 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_1_3 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_1_3 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_1_3 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_1_3 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_1_3 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_1_3 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_1_3 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_1_3 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_1_3 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_1_3 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_1_3 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_1_3 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_1_3 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_1_3 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_1_3 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_1_3 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_1_3 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_1_3 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_1_3 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_1_3 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_1_3 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_1_3 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_1_3 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_1_3 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_1_3 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_1_3 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_1_3 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_1_3 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_1_3 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_1_3 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_1_3 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_1_3 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_1_3 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_1_3 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_1_3 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_1_3 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_1_3 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_1_3 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_1_3 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_1_3 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_1_3 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_1_3 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_1_3 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_1_3 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_1_3 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_1_3 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_1_3 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_1_3 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_1_3 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_1_3 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_1_3 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_1_3 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_1_3 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_1_3 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_1_3 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_1_3 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_1_3 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_1_3 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_1_3 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_1_3 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_1_3 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_1_3 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_1_3 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_1_3 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_1_3 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_1_3 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_1_3 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_1_3 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_1_3 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_1_3 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_1_3 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_1_3 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_1_3 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_1_3 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_1_3 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_1_3 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_1_3 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_1_3 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_1_3 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_1_3 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_1_3 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_1_3 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_1_3 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_1_3 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_1_3 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_1_3 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_1_3 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_1_3 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_1_3 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_1_3 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_1_3 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_1_3 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_1_3 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_1_3 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_1_3 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_1_3 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_1_3 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_1_3 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_1_3 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_1_3 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_1_3 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_1_3 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_1_3 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_1_3 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_1_3 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_1_3 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_1_3 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_1_3 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_1_3 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_1_3 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_1_3 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_1_3 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_1_3 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_1_3 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_1_3 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_1_3 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_1_3 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_1_3 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_1_3 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_1_3 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_1_3 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_1_3 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_1_3 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_1_3 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_1_3 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_1_3 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_1_3 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_1_3 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_1_3 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_1_3 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_1_3 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_1_3 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_1_3 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_1_3 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_1_3 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_1_3 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_1_3 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_1_3 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_1_3 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_1_3 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_1_3 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_1_3 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_1_3 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_1_3 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_1_3 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_1_3 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_1_3 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_1_3 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_1_3 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_1_3 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_1_3 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_1_3 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_1_3 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_1_3 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_1_3 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_1_3 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_1_3 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_1_3 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_1_3 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_1_3 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_1_3 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_1_3 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_1_3 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_1_3 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_1_3 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_1_3 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_1_3 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_1_3 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_1_3 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_1_3 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_1_3 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_1_3 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_1_3 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_1_3 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_1_3 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_1_3 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_1_3 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_1_3 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_1_3 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_1_3 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_1_3 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_1_3 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_1_3 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_1_3 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_1_3 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_1_3 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_1_3 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_1_3 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_1_3 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_1_3 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_1_3 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_1_3 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_1_3 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_1_3 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_1_3 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_1_3 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_1_3 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_1_3 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_1_3 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_1_3 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_1_3 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_1_3 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_1_3 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_1_3 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_1_3 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_1_3 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_1_3 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_1_3 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_1_3 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_1_3 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_1_3 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_1_3 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_1_3 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_1_3 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_1_3 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_1_3 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_1_3 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_1_3 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_1_3 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_1_3 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_1_3 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_1_3 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_1_3 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_1_3 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_1_3 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_1_3 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_1_3 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_12_1 <= out0_124(12);

  
  s_12 <= sbox(0) WHEN out0_12_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_12_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_12_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_12_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_12_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_12_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_12_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_12_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_12_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_12_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_12_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_12_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_12_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_12_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_12_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_12_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_12_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_12_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_12_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_12_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_12_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_12_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_12_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_12_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_12_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_12_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_12_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_12_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_12_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_12_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_12_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_12_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_12_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_12_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_12_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_12_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_12_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_12_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_12_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_12_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_12_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_12_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_12_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_12_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_12_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_12_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_12_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_12_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_12_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_12_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_12_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_12_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_12_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_12_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_12_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_12_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_12_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_12_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_12_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_12_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_12_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_12_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_12_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_12_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_12_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_12_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_12_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_12_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_12_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_12_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_12_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_12_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_12_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_12_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_12_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_12_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_12_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_12_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_12_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_12_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_12_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_12_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_12_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_12_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_12_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_12_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_12_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_12_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_12_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_12_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_12_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_12_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_12_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_12_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_12_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_12_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_12_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_12_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_12_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_12_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_12_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_12_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_12_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_12_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_12_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_12_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_12_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_12_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_12_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_12_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_12_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_12_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_12_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_12_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_12_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_12_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_12_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_12_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_12_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_12_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_12_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_12_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_12_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_12_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_12_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_12_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_12_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_12_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_12_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_12_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_12_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_12_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_12_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_12_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_12_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_12_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_12_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_12_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_12_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_12_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_12_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_12_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_12_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_12_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_12_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_12_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_12_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_12_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_12_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_12_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_12_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_12_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_12_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_12_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_12_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_12_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_12_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_12_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_12_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_12_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_12_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_12_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_12_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_12_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_12_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_12_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_12_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_12_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_12_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_12_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_12_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_12_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_12_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_12_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_12_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_12_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_12_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_12_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_12_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_12_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_12_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_12_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_12_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_12_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_12_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_12_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_12_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_12_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_12_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_12_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_12_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_12_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_12_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_12_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_12_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_12_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_12_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_12_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_12_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_12_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_12_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_12_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_12_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_12_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_12_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_12_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_12_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_12_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_12_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_12_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_12_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_12_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_12_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_12_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_12_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_12_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_12_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_12_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_12_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_12_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_12_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_12_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_12_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_12_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_12_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_12_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_12_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_12_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_12_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_12_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_12_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_12_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_12_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_12_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_12_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_12_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_12_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_12_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_12_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_12_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_12_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_12_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_12_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_12_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_12_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_12_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_12_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_12_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_12_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_12_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_12_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_12_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_12_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_12_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_12_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_7_1 <= out0_124(7);

  
  s_7 <= sbox(0) WHEN out0_7_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_7_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_7_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_7_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_7_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_7_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_7_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_7_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_7_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_7_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_7_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_7_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_7_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_7_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_7_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_7_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_7_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_7_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_7_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_7_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_7_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_7_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_7_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_7_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_7_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_7_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_7_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_7_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_7_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_7_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_7_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_7_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_7_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_7_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_7_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_7_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_7_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_7_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_7_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_7_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_7_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_7_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_7_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_7_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_7_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_7_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_7_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_7_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_7_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_7_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_7_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_7_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_7_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_7_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_7_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_7_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_7_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_7_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_7_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_7_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_7_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_7_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_7_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_7_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_7_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_7_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_7_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_7_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_7_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_7_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_7_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_7_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_7_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_7_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_7_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_7_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_7_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_7_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_7_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_7_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_7_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_7_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_7_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_7_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_7_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_7_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_7_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_7_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_7_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_7_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_7_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_7_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_7_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_7_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_7_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_7_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_7_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_7_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_7_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_7_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_7_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_7_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_7_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_7_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_7_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_7_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_7_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_7_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_7_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_7_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_7_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_7_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_7_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_7_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_7_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_7_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_7_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_7_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_7_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_7_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_7_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_7_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_7_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_7_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_7_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_7_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_7_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_7_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_7_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_7_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_7_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_7_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_7_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_7_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_7_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_7_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_7_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_7_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_7_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_7_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_7_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_7_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_7_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_7_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_7_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_7_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_7_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_7_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_7_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_7_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_7_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_7_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_7_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_7_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_7_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_7_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_7_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_7_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_7_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_7_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_7_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_7_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_7_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_7_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_7_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_7_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_7_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_7_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_7_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_7_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_7_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_7_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_7_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_7_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_7_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_7_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_7_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_7_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_7_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_7_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_7_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_7_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_7_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_7_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_7_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_7_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_7_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_7_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_7_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_7_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_7_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_7_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_7_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_7_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_7_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_7_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_7_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_7_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_7_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_7_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_7_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_7_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_7_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_7_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_7_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_7_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_7_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_7_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_7_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_7_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_7_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_7_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_7_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_7_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_7_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_7_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_7_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_7_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_7_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_7_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_7_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_7_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_7_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_7_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_7_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_7_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_7_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_7_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_7_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_7_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_7_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_7_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_7_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_7_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_7_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_7_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_7_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_7_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_7_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_7_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_7_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_7_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_7_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_7_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_7_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_7_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_7_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_7_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_7_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_7_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_7_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_7_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_7_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_7_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_7_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_2_3 <= out0_124(2);

  
  s_2 <= sbox(0) WHEN out0_2_3 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_2_3 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_2_3 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_2_3 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_2_3 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_2_3 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_2_3 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_2_3 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_2_3 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_2_3 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_2_3 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_2_3 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_2_3 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_2_3 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_2_3 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_2_3 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_2_3 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_2_3 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_2_3 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_2_3 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_2_3 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_2_3 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_2_3 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_2_3 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_2_3 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_2_3 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_2_3 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_2_3 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_2_3 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_2_3 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_2_3 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_2_3 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_2_3 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_2_3 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_2_3 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_2_3 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_2_3 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_2_3 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_2_3 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_2_3 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_2_3 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_2_3 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_2_3 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_2_3 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_2_3 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_2_3 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_2_3 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_2_3 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_2_3 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_2_3 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_2_3 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_2_3 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_2_3 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_2_3 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_2_3 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_2_3 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_2_3 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_2_3 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_2_3 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_2_3 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_2_3 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_2_3 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_2_3 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_2_3 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_2_3 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_2_3 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_2_3 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_2_3 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_2_3 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_2_3 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_2_3 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_2_3 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_2_3 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_2_3 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_2_3 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_2_3 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_2_3 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_2_3 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_2_3 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_2_3 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_2_3 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_2_3 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_2_3 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_2_3 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_2_3 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_2_3 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_2_3 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_2_3 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_2_3 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_2_3 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_2_3 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_2_3 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_2_3 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_2_3 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_2_3 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_2_3 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_2_3 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_2_3 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_2_3 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_2_3 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_2_3 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_2_3 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_2_3 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_2_3 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_2_3 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_2_3 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_2_3 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_2_3 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_2_3 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_2_3 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_2_3 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_2_3 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_2_3 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_2_3 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_2_3 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_2_3 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_2_3 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_2_3 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_2_3 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_2_3 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_2_3 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_2_3 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_2_3 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_2_3 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_2_3 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_2_3 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_2_3 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_2_3 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_2_3 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_2_3 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_2_3 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_2_3 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_2_3 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_2_3 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_2_3 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_2_3 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_2_3 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_2_3 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_2_3 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_2_3 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_2_3 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_2_3 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_2_3 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_2_3 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_2_3 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_2_3 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_2_3 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_2_3 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_2_3 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_2_3 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_2_3 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_2_3 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_2_3 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_2_3 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_2_3 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_2_3 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_2_3 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_2_3 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_2_3 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_2_3 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_2_3 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_2_3 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_2_3 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_2_3 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_2_3 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_2_3 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_2_3 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_2_3 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_2_3 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_2_3 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_2_3 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_2_3 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_2_3 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_2_3 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_2_3 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_2_3 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_2_3 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_2_3 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_2_3 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_2_3 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_2_3 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_2_3 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_2_3 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_2_3 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_2_3 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_2_3 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_2_3 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_2_3 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_2_3 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_2_3 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_2_3 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_2_3 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_2_3 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_2_3 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_2_3 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_2_3 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_2_3 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_2_3 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_2_3 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_2_3 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_2_3 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_2_3 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_2_3 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_2_3 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_2_3 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_2_3 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_2_3 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_2_3 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_2_3 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_2_3 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_2_3 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_2_3 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_2_3 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_2_3 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_2_3 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_2_3 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_2_3 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_2_3 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_2_3 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_2_3 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_2_3 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_2_3 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_2_3 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_2_3 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_2_3 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_2_3 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_2_3 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_2_3 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_2_3 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_2_3 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_2_3 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_2_3 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_2_3 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_2_3 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_2_3 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_2_3 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_2_3 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_2_3 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_2_3 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_2_3 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_2_3 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_2_3 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_2_3 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_2_3 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_2_3 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_2_3 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_2_3 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_2_3 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_2_3 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_2_3 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_2_3 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_2_3 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_2_3 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_2_3 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_2_3 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_13_1 <= out0_124(13);

  
  s_13 <= sbox(0) WHEN out0_13_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_13_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_13_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_13_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_13_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_13_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_13_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_13_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_13_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_13_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_13_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_13_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_13_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_13_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_13_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_13_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_13_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_13_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_13_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_13_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_13_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_13_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_13_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_13_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_13_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_13_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_13_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_13_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_13_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_13_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_13_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_13_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_13_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_13_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_13_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_13_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_13_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_13_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_13_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_13_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_13_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_13_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_13_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_13_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_13_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_13_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_13_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_13_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_13_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_13_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_13_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_13_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_13_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_13_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_13_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_13_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_13_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_13_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_13_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_13_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_13_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_13_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_13_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_13_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_13_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_13_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_13_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_13_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_13_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_13_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_13_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_13_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_13_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_13_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_13_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_13_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_13_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_13_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_13_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_13_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_13_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_13_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_13_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_13_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_13_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_13_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_13_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_13_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_13_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_13_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_13_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_13_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_13_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_13_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_13_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_13_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_13_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_13_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_13_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_13_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_13_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_13_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_13_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_13_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_13_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_13_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_13_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_13_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_13_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_13_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_13_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_13_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_13_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_13_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_13_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_13_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_13_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_13_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_13_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_13_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_13_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_13_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_13_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_13_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_13_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_13_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_13_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_13_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_13_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_13_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_13_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_13_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_13_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_13_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_13_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_13_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_13_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_13_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_13_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_13_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_13_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_13_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_13_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_13_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_13_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_13_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_13_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_13_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_13_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_13_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_13_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_13_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_13_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_13_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_13_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_13_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_13_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_13_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_13_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_13_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_13_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_13_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_13_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_13_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_13_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_13_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_13_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_13_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_13_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_13_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_13_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_13_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_13_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_13_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_13_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_13_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_13_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_13_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_13_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_13_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_13_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_13_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_13_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_13_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_13_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_13_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_13_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_13_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_13_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_13_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_13_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_13_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_13_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_13_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_13_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_13_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_13_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_13_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_13_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_13_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_13_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_13_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_13_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_13_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_13_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_13_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_13_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_13_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_13_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_13_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_13_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_13_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_13_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_13_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_13_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_13_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_13_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_13_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_13_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_13_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_13_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_13_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_13_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_13_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_13_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_13_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_13_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_13_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_13_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_13_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_13_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_13_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_13_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_13_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_13_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_13_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_13_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_13_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_13_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_13_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_13_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_13_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_13_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_13_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_13_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_13_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_13_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_13_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_13_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_13_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_13_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_13_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_13_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_13_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_13_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_8_1 <= out0_124(8);

  
  s_8 <= sbox(0) WHEN out0_8_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_8_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_8_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_8_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_8_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_8_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_8_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_8_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_8_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_8_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_8_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_8_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_8_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_8_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_8_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_8_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_8_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_8_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_8_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_8_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_8_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_8_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_8_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_8_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_8_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_8_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_8_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_8_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_8_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_8_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_8_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_8_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_8_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_8_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_8_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_8_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_8_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_8_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_8_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_8_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_8_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_8_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_8_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_8_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_8_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_8_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_8_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_8_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_8_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_8_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_8_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_8_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_8_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_8_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_8_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_8_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_8_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_8_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_8_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_8_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_8_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_8_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_8_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_8_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_8_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_8_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_8_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_8_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_8_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_8_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_8_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_8_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_8_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_8_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_8_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_8_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_8_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_8_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_8_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_8_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_8_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_8_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_8_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_8_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_8_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_8_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_8_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_8_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_8_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_8_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_8_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_8_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_8_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_8_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_8_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_8_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_8_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_8_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_8_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_8_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_8_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_8_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_8_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_8_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_8_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_8_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_8_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_8_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_8_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_8_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_8_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_8_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_8_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_8_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_8_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_8_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_8_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_8_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_8_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_8_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_8_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_8_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_8_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_8_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_8_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_8_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_8_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_8_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_8_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_8_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_8_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_8_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_8_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_8_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_8_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_8_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_8_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_8_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_8_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_8_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_8_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_8_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_8_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_8_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_8_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_8_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_8_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_8_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_8_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_8_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_8_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_8_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_8_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_8_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_8_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_8_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_8_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_8_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_8_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_8_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_8_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_8_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_8_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_8_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_8_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_8_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_8_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_8_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_8_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_8_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_8_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_8_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_8_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_8_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_8_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_8_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_8_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_8_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_8_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_8_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_8_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_8_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_8_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_8_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_8_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_8_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_8_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_8_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_8_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_8_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_8_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_8_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_8_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_8_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_8_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_8_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_8_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_8_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_8_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_8_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_8_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_8_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_8_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_8_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_8_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_8_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_8_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_8_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_8_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_8_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_8_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_8_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_8_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_8_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_8_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_8_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_8_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_8_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_8_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_8_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_8_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_8_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_8_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_8_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_8_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_8_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_8_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_8_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_8_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_8_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_8_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_8_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_8_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_8_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_8_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_8_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_8_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_8_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_8_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_8_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_8_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_8_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_8_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_8_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_8_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_8_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_8_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_8_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_8_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_8_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_8_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_8_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_8_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_8_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_8_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_3_3 <= out0_124(3);

  
  s_3 <= sbox(0) WHEN out0_3_3 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_3_3 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_3_3 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_3_3 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_3_3 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_3_3 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_3_3 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_3_3 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_3_3 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_3_3 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_3_3 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_3_3 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_3_3 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_3_3 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_3_3 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_3_3 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_3_3 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_3_3 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_3_3 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_3_3 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_3_3 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_3_3 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_3_3 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_3_3 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_3_3 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_3_3 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_3_3 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_3_3 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_3_3 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_3_3 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_3_3 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_3_3 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_3_3 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_3_3 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_3_3 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_3_3 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_3_3 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_3_3 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_3_3 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_3_3 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_3_3 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_3_3 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_3_3 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_3_3 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_3_3 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_3_3 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_3_3 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_3_3 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_3_3 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_3_3 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_3_3 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_3_3 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_3_3 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_3_3 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_3_3 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_3_3 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_3_3 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_3_3 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_3_3 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_3_3 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_3_3 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_3_3 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_3_3 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_3_3 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_3_3 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_3_3 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_3_3 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_3_3 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_3_3 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_3_3 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_3_3 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_3_3 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_3_3 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_3_3 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_3_3 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_3_3 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_3_3 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_3_3 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_3_3 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_3_3 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_3_3 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_3_3 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_3_3 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_3_3 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_3_3 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_3_3 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_3_3 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_3_3 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_3_3 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_3_3 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_3_3 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_3_3 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_3_3 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_3_3 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_3_3 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_3_3 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_3_3 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_3_3 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_3_3 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_3_3 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_3_3 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_3_3 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_3_3 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_3_3 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_3_3 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_3_3 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_3_3 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_3_3 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_3_3 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_3_3 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_3_3 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_3_3 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_3_3 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_3_3 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_3_3 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_3_3 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_3_3 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_3_3 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_3_3 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_3_3 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_3_3 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_3_3 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_3_3 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_3_3 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_3_3 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_3_3 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_3_3 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_3_3 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_3_3 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_3_3 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_3_3 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_3_3 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_3_3 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_3_3 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_3_3 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_3_3 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_3_3 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_3_3 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_3_3 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_3_3 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_3_3 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_3_3 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_3_3 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_3_3 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_3_3 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_3_3 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_3_3 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_3_3 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_3_3 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_3_3 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_3_3 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_3_3 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_3_3 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_3_3 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_3_3 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_3_3 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_3_3 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_3_3 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_3_3 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_3_3 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_3_3 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_3_3 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_3_3 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_3_3 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_3_3 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_3_3 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_3_3 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_3_3 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_3_3 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_3_3 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_3_3 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_3_3 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_3_3 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_3_3 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_3_3 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_3_3 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_3_3 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_3_3 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_3_3 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_3_3 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_3_3 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_3_3 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_3_3 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_3_3 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_3_3 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_3_3 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_3_3 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_3_3 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_3_3 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_3_3 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_3_3 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_3_3 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_3_3 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_3_3 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_3_3 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_3_3 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_3_3 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_3_3 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_3_3 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_3_3 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_3_3 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_3_3 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_3_3 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_3_3 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_3_3 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_3_3 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_3_3 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_3_3 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_3_3 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_3_3 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_3_3 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_3_3 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_3_3 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_3_3 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_3_3 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_3_3 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_3_3 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_3_3 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_3_3 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_3_3 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_3_3 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_3_3 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_3_3 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_3_3 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_3_3 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_3_3 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_3_3 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_3_3 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_3_3 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_3_3 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_3_3 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_3_3 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_3_3 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_3_3 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_3_3 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_3_3 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_3_3 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_3_3 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_3_3 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_3_3 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_3_3 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_3_3 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_3_3 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_3_3 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_3_3 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_3_3 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_3_3 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_3_3 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_3_3 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_3_3 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_3_3 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_3_3 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_3_3 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_3_3 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_3_3 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_14_1 <= out0_124(14);

  
  s_14 <= sbox(0) WHEN out0_14_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_14_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_14_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_14_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_14_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_14_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_14_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_14_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_14_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_14_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_14_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_14_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_14_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_14_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_14_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_14_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_14_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_14_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_14_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_14_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_14_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_14_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_14_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_14_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_14_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_14_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_14_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_14_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_14_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_14_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_14_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_14_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_14_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_14_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_14_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_14_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_14_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_14_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_14_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_14_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_14_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_14_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_14_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_14_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_14_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_14_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_14_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_14_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_14_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_14_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_14_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_14_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_14_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_14_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_14_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_14_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_14_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_14_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_14_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_14_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_14_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_14_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_14_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_14_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_14_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_14_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_14_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_14_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_14_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_14_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_14_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_14_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_14_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_14_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_14_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_14_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_14_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_14_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_14_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_14_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_14_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_14_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_14_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_14_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_14_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_14_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_14_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_14_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_14_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_14_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_14_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_14_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_14_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_14_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_14_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_14_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_14_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_14_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_14_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_14_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_14_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_14_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_14_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_14_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_14_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_14_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_14_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_14_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_14_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_14_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_14_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_14_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_14_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_14_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_14_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_14_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_14_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_14_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_14_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_14_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_14_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_14_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_14_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_14_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_14_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_14_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_14_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_14_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_14_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_14_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_14_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_14_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_14_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_14_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_14_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_14_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_14_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_14_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_14_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_14_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_14_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_14_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_14_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_14_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_14_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_14_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_14_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_14_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_14_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_14_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_14_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_14_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_14_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_14_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_14_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_14_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_14_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_14_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_14_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_14_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_14_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_14_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_14_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_14_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_14_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_14_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_14_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_14_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_14_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_14_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_14_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_14_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_14_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_14_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_14_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_14_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_14_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_14_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_14_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_14_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_14_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_14_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_14_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_14_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_14_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_14_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_14_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_14_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_14_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_14_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_14_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_14_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_14_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_14_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_14_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_14_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_14_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_14_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_14_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_14_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_14_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_14_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_14_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_14_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_14_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_14_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_14_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_14_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_14_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_14_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_14_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_14_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_14_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_14_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_14_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_14_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_14_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_14_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_14_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_14_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_14_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_14_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_14_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_14_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_14_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_14_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_14_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_14_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_14_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_14_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_14_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_14_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_14_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_14_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_14_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_14_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_14_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_14_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_14_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_14_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_14_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_14_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_14_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_14_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_14_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_14_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_14_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_14_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_14_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_14_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_14_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_14_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_14_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_14_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_14_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_9_1 <= out0_124(9);

  
  s_9 <= sbox(0) WHEN out0_9_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_9_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_9_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_9_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_9_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_9_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_9_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_9_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_9_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_9_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_9_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_9_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_9_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_9_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_9_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_9_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_9_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_9_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_9_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_9_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_9_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_9_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_9_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_9_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_9_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_9_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_9_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_9_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_9_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_9_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_9_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_9_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_9_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_9_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_9_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_9_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_9_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_9_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_9_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_9_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_9_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_9_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_9_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_9_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_9_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_9_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_9_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_9_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_9_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_9_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_9_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_9_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_9_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_9_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_9_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_9_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_9_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_9_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_9_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_9_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_9_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_9_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_9_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_9_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_9_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_9_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_9_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_9_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_9_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_9_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_9_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_9_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_9_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_9_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_9_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_9_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_9_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_9_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_9_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_9_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_9_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_9_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_9_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_9_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_9_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_9_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_9_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_9_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_9_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_9_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_9_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_9_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_9_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_9_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_9_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_9_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_9_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_9_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_9_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_9_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_9_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_9_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_9_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_9_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_9_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_9_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_9_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_9_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_9_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_9_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_9_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_9_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_9_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_9_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_9_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_9_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_9_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_9_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_9_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_9_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_9_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_9_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_9_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_9_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_9_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_9_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_9_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_9_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_9_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_9_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_9_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_9_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_9_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_9_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_9_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_9_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_9_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_9_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_9_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_9_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_9_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_9_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_9_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_9_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_9_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_9_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_9_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_9_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_9_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_9_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_9_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_9_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_9_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_9_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_9_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_9_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_9_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_9_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_9_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_9_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_9_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_9_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_9_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_9_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_9_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_9_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_9_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_9_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_9_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_9_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_9_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_9_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_9_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_9_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_9_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_9_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_9_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_9_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_9_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_9_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_9_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_9_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_9_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_9_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_9_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_9_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_9_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_9_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_9_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_9_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_9_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_9_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_9_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_9_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_9_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_9_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_9_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_9_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_9_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_9_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_9_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_9_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_9_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_9_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_9_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_9_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_9_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_9_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_9_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_9_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_9_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_9_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_9_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_9_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_9_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_9_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_9_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_9_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_9_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_9_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_9_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_9_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_9_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_9_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_9_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_9_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_9_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_9_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_9_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_9_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_9_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_9_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_9_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_9_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_9_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_9_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_9_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_9_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_9_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_9_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_9_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_9_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_9_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_9_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_9_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_9_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_9_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_9_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_9_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_9_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_9_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_9_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_9_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_9_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_9_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_4_1 <= out0_124(4);

  
  s_4 <= sbox(0) WHEN out0_4_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_4_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_4_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_4_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_4_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_4_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_4_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_4_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_4_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_4_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_4_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_4_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_4_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_4_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_4_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_4_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_4_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_4_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_4_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_4_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_4_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_4_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_4_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_4_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_4_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_4_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_4_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_4_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_4_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_4_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_4_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_4_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_4_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_4_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_4_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_4_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_4_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_4_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_4_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_4_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_4_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_4_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_4_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_4_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_4_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_4_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_4_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_4_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_4_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_4_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_4_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_4_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_4_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_4_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_4_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_4_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_4_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_4_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_4_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_4_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_4_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_4_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_4_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_4_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_4_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_4_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_4_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_4_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_4_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_4_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_4_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_4_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_4_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_4_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_4_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_4_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_4_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_4_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_4_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_4_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_4_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_4_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_4_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_4_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_4_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_4_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_4_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_4_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_4_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_4_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_4_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_4_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_4_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_4_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_4_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_4_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_4_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_4_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_4_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_4_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_4_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_4_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_4_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_4_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_4_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_4_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_4_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_4_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_4_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_4_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_4_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_4_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_4_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_4_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_4_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_4_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_4_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_4_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_4_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_4_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_4_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_4_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_4_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_4_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_4_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_4_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_4_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_4_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_4_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_4_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_4_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_4_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_4_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_4_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_4_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_4_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_4_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_4_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_4_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_4_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_4_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_4_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_4_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_4_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_4_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_4_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_4_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_4_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_4_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_4_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_4_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_4_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_4_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_4_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_4_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_4_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_4_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_4_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_4_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_4_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_4_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_4_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_4_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_4_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_4_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_4_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_4_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_4_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_4_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_4_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_4_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_4_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_4_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_4_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_4_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_4_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_4_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_4_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_4_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_4_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_4_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_4_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_4_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_4_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_4_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_4_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_4_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_4_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_4_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_4_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_4_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_4_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_4_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_4_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_4_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_4_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_4_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_4_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_4_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_4_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_4_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_4_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_4_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_4_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_4_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_4_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_4_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_4_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_4_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_4_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_4_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_4_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_4_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_4_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_4_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_4_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_4_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_4_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_4_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_4_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_4_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_4_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_4_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_4_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_4_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_4_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_4_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_4_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_4_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_4_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_4_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_4_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_4_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_4_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_4_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_4_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_4_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_4_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_4_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_4_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_4_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_4_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_4_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_4_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_4_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_4_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_4_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_4_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_4_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_4_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_4_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_4_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_4_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_4_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_4_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_15_1 <= out0_124(15);

  
  s_15 <= sbox(0) WHEN out0_15_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_15_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_15_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_15_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_15_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_15_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_15_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_15_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_15_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_15_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_15_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_15_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_15_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_15_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_15_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_15_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_15_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_15_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_15_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_15_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_15_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_15_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_15_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_15_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_15_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_15_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_15_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_15_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_15_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_15_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_15_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_15_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_15_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_15_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_15_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_15_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_15_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_15_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_15_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_15_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_15_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_15_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_15_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_15_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_15_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_15_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_15_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_15_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_15_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_15_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_15_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_15_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_15_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_15_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_15_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_15_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_15_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_15_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_15_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_15_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_15_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_15_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_15_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_15_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_15_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_15_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_15_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_15_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_15_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_15_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_15_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_15_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_15_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_15_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_15_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_15_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_15_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_15_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_15_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_15_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_15_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_15_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_15_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_15_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_15_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_15_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_15_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_15_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_15_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_15_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_15_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_15_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_15_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_15_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_15_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_15_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_15_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_15_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_15_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_15_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_15_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_15_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_15_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_15_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_15_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_15_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_15_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_15_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_15_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_15_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_15_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_15_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_15_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_15_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_15_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_15_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_15_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_15_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_15_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_15_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_15_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_15_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_15_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_15_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_15_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_15_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_15_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_15_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_15_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_15_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_15_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_15_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_15_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_15_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_15_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_15_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_15_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_15_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_15_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_15_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_15_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_15_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_15_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_15_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_15_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_15_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_15_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_15_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_15_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_15_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_15_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_15_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_15_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_15_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_15_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_15_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_15_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_15_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_15_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_15_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_15_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_15_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_15_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_15_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_15_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_15_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_15_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_15_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_15_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_15_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_15_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_15_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_15_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_15_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_15_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_15_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_15_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_15_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_15_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_15_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_15_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_15_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_15_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_15_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_15_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_15_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_15_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_15_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_15_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_15_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_15_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_15_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_15_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_15_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_15_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_15_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_15_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_15_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_15_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_15_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_15_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_15_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_15_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_15_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_15_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_15_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_15_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_15_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_15_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_15_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_15_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_15_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_15_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_15_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_15_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_15_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_15_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_15_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_15_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_15_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_15_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_15_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_15_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_15_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_15_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_15_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_15_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_15_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_15_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_15_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_15_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_15_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_15_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_15_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_15_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_15_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_15_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_15_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_15_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_15_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_15_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_15_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_15_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_15_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_15_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_15_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_15_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_15_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_15_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_15_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_15_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_15_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_15_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_15_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_15_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_10_1 <= out0_124(10);

  
  s_10 <= sbox(0) WHEN out0_10_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_10_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_10_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_10_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_10_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_10_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_10_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_10_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_10_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_10_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_10_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_10_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_10_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_10_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_10_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_10_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_10_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_10_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_10_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_10_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_10_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_10_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_10_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_10_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_10_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_10_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_10_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_10_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_10_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_10_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_10_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_10_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_10_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_10_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_10_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_10_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_10_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_10_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_10_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_10_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_10_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_10_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_10_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_10_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_10_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_10_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_10_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_10_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_10_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_10_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_10_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_10_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_10_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_10_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_10_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_10_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_10_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_10_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_10_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_10_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_10_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_10_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_10_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_10_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_10_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_10_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_10_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_10_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_10_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_10_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_10_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_10_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_10_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_10_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_10_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_10_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_10_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_10_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_10_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_10_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_10_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_10_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_10_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_10_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_10_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_10_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_10_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_10_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_10_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_10_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_10_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_10_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_10_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_10_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_10_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_10_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_10_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_10_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_10_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_10_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_10_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_10_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_10_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_10_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_10_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_10_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_10_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_10_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_10_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_10_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_10_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_10_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_10_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_10_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_10_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_10_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_10_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_10_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_10_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_10_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_10_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_10_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_10_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_10_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_10_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_10_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_10_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_10_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_10_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_10_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_10_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_10_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_10_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_10_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_10_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_10_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_10_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_10_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_10_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_10_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_10_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_10_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_10_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_10_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_10_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_10_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_10_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_10_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_10_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_10_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_10_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_10_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_10_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_10_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_10_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_10_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_10_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_10_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_10_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_10_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_10_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_10_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_10_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_10_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_10_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_10_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_10_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_10_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_10_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_10_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_10_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_10_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_10_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_10_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_10_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_10_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_10_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_10_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_10_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_10_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_10_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_10_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_10_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_10_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_10_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_10_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_10_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_10_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_10_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_10_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_10_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_10_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_10_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_10_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_10_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_10_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_10_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_10_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_10_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_10_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_10_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_10_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_10_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_10_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_10_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_10_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_10_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_10_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_10_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_10_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_10_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_10_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_10_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_10_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_10_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_10_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_10_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_10_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_10_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_10_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_10_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_10_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_10_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_10_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_10_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_10_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_10_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_10_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_10_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_10_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_10_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_10_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_10_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_10_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_10_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_10_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_10_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_10_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_10_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_10_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_10_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_10_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_10_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_10_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_10_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_10_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_10_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_10_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_10_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_10_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_10_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_10_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_10_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_10_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_10_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_5_1 <= out0_124(5);

  
  s_5 <= sbox(0) WHEN out0_5_1 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_5_1 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_5_1 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_5_1 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_5_1 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_5_1 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_5_1 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_5_1 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_5_1 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_5_1 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_5_1 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_5_1 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_5_1 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_5_1 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_5_1 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_5_1 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_5_1 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_5_1 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_5_1 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_5_1 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_5_1 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_5_1 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_5_1 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_5_1 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_5_1 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_5_1 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_5_1 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_5_1 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_5_1 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_5_1 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_5_1 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_5_1 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_5_1 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_5_1 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_5_1 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_5_1 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_5_1 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_5_1 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_5_1 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_5_1 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_5_1 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_5_1 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_5_1 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_5_1 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_5_1 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_5_1 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_5_1 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_5_1 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_5_1 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_5_1 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_5_1 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_5_1 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_5_1 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_5_1 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_5_1 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_5_1 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_5_1 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_5_1 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_5_1 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_5_1 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_5_1 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_5_1 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_5_1 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_5_1 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_5_1 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_5_1 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_5_1 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_5_1 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_5_1 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_5_1 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_5_1 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_5_1 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_5_1 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_5_1 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_5_1 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_5_1 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_5_1 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_5_1 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_5_1 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_5_1 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_5_1 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_5_1 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_5_1 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_5_1 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_5_1 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_5_1 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_5_1 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_5_1 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_5_1 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_5_1 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_5_1 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_5_1 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_5_1 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_5_1 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_5_1 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_5_1 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_5_1 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_5_1 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_5_1 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_5_1 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_5_1 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_5_1 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_5_1 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_5_1 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_5_1 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_5_1 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_5_1 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_5_1 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_5_1 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_5_1 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_5_1 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_5_1 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_5_1 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_5_1 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_5_1 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_5_1 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_5_1 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_5_1 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_5_1 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_5_1 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_5_1 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_5_1 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_5_1 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_5_1 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_5_1 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_5_1 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_5_1 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_5_1 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_5_1 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_5_1 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_5_1 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_5_1 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_5_1 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_5_1 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_5_1 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_5_1 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_5_1 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_5_1 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_5_1 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_5_1 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_5_1 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_5_1 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_5_1 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_5_1 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_5_1 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_5_1 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_5_1 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_5_1 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_5_1 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_5_1 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_5_1 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_5_1 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_5_1 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_5_1 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_5_1 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_5_1 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_5_1 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_5_1 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_5_1 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_5_1 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_5_1 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_5_1 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_5_1 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_5_1 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_5_1 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_5_1 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_5_1 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_5_1 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_5_1 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_5_1 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_5_1 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_5_1 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_5_1 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_5_1 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_5_1 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_5_1 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_5_1 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_5_1 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_5_1 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_5_1 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_5_1 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_5_1 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_5_1 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_5_1 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_5_1 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_5_1 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_5_1 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_5_1 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_5_1 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_5_1 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_5_1 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_5_1 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_5_1 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_5_1 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_5_1 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_5_1 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_5_1 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_5_1 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_5_1 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_5_1 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_5_1 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_5_1 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_5_1 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_5_1 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_5_1 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_5_1 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_5_1 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_5_1 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_5_1 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_5_1 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_5_1 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_5_1 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_5_1 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_5_1 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_5_1 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_5_1 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_5_1 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_5_1 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_5_1 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_5_1 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_5_1 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_5_1 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_5_1 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_5_1 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_5_1 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_5_1 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_5_1 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_5_1 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_5_1 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_5_1 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_5_1 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_5_1 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_5_1 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_5_1 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_5_1 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_5_1 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_5_1 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_5_1 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_5_1 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_5_1 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_5_1 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_5_1 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_5_1 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_5_1 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_5_1 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_5_1 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_5_1 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_5_1 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_5_1 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_5_1 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_5_1 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_5_1 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_5_1 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_5_1 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_5_1 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  out0_125(0) <= s_s_1(0);
  out0_125(1) <= s_s_1(1);
  out0_125(2) <= s_s_1(2);
  out0_125(3) <= s_s_1(3);
  out0_125(4) <= s_s_1(4);
  out0_125(5) <= s_s_1(5);
  out0_125(6) <= s_s_1(6);
  out0_125(7) <= s_s_1(7);
  out0_125(8) <= s_s_1(8);
  out0_125(9) <= s_s_1(9);
  out0_125(10) <= s_s_1(10);
  out0_125(11) <= s_s_1(11);
  out0_125(12) <= s_s_1(12);
  out0_125(13) <= s_s_1(13);
  out0_125(14) <= s_s_1(14);
  out0_125(15) <= s_s_1(15);

  out0_126(0) <= resize(out0_125(0), 16);
  out0_126(1) <= resize(out0_125(1), 16);
  out0_126(2) <= resize(out0_125(2), 16);
  out0_126(3) <= resize(out0_125(3), 16);
  out0_126(4) <= resize(out0_125(4), 16);
  out0_126(5) <= resize(out0_125(5), 16);
  out0_126(6) <= resize(out0_125(6), 16);
  out0_126(7) <= resize(out0_125(7), 16);
  out0_126(8) <= resize(out0_125(8), 16);
  out0_126(9) <= resize(out0_125(9), 16);
  out0_126(10) <= resize(out0_125(10), 16);
  out0_126(11) <= resize(out0_125(11), 16);
  out0_126(12) <= resize(out0_125(12), 16);
  out0_126(13) <= resize(out0_125(13), 16);
  out0_126(14) <= resize(out0_125(14), 16);
  out0_126(15) <= resize(out0_125(15), 16);

  out0_124(0) <= out0_126(0) + const_expression_26;
  out0_124(1) <= out0_126(1) + const_expression_26;
  out0_124(2) <= out0_126(2) + const_expression_26;
  out0_124(3) <= out0_126(3) + const_expression_26;
  out0_124(4) <= out0_126(4) + const_expression_26;
  out0_124(5) <= out0_126(5) + const_expression_26;
  out0_124(6) <= out0_126(6) + const_expression_26;
  out0_124(7) <= out0_126(7) + const_expression_26;
  out0_124(8) <= out0_126(8) + const_expression_26;
  out0_124(9) <= out0_126(9) + const_expression_26;
  out0_124(10) <= out0_126(10) + const_expression_26;
  out0_124(11) <= out0_126(11) + const_expression_26;
  out0_124(12) <= out0_126(12) + const_expression_26;
  out0_124(13) <= out0_126(13) + const_expression_26;
  out0_124(14) <= out0_126(14) + const_expression_26;
  out0_124(15) <= out0_126(15) + const_expression_26;

  out0_0_2 <= out0_124(0);

  
  s_0 <= sbox(0) WHEN out0_0_2 = to_unsigned(16#0001#, 16) ELSE
      sbox(1) WHEN out0_0_2 = to_unsigned(16#0002#, 16) ELSE
      sbox(2) WHEN out0_0_2 = to_unsigned(16#0003#, 16) ELSE
      sbox(3) WHEN out0_0_2 = to_unsigned(16#0004#, 16) ELSE
      sbox(4) WHEN out0_0_2 = to_unsigned(16#0005#, 16) ELSE
      sbox(5) WHEN out0_0_2 = to_unsigned(16#0006#, 16) ELSE
      sbox(6) WHEN out0_0_2 = to_unsigned(16#0007#, 16) ELSE
      sbox(7) WHEN out0_0_2 = to_unsigned(16#0008#, 16) ELSE
      sbox(8) WHEN out0_0_2 = to_unsigned(16#0009#, 16) ELSE
      sbox(9) WHEN out0_0_2 = to_unsigned(16#000A#, 16) ELSE
      sbox(10) WHEN out0_0_2 = to_unsigned(16#000B#, 16) ELSE
      sbox(11) WHEN out0_0_2 = to_unsigned(16#000C#, 16) ELSE
      sbox(12) WHEN out0_0_2 = to_unsigned(16#000D#, 16) ELSE
      sbox(13) WHEN out0_0_2 = to_unsigned(16#000E#, 16) ELSE
      sbox(14) WHEN out0_0_2 = to_unsigned(16#000F#, 16) ELSE
      sbox(15) WHEN out0_0_2 = to_unsigned(16#0010#, 16) ELSE
      sbox(16) WHEN out0_0_2 = to_unsigned(16#0011#, 16) ELSE
      sbox(17) WHEN out0_0_2 = to_unsigned(16#0012#, 16) ELSE
      sbox(18) WHEN out0_0_2 = to_unsigned(16#0013#, 16) ELSE
      sbox(19) WHEN out0_0_2 = to_unsigned(16#0014#, 16) ELSE
      sbox(20) WHEN out0_0_2 = to_unsigned(16#0015#, 16) ELSE
      sbox(21) WHEN out0_0_2 = to_unsigned(16#0016#, 16) ELSE
      sbox(22) WHEN out0_0_2 = to_unsigned(16#0017#, 16) ELSE
      sbox(23) WHEN out0_0_2 = to_unsigned(16#0018#, 16) ELSE
      sbox(24) WHEN out0_0_2 = to_unsigned(16#0019#, 16) ELSE
      sbox(25) WHEN out0_0_2 = to_unsigned(16#001A#, 16) ELSE
      sbox(26) WHEN out0_0_2 = to_unsigned(16#001B#, 16) ELSE
      sbox(27) WHEN out0_0_2 = to_unsigned(16#001C#, 16) ELSE
      sbox(28) WHEN out0_0_2 = to_unsigned(16#001D#, 16) ELSE
      sbox(29) WHEN out0_0_2 = to_unsigned(16#001E#, 16) ELSE
      sbox(30) WHEN out0_0_2 = to_unsigned(16#001F#, 16) ELSE
      sbox(31) WHEN out0_0_2 = to_unsigned(16#0020#, 16) ELSE
      sbox(32) WHEN out0_0_2 = to_unsigned(16#0021#, 16) ELSE
      sbox(33) WHEN out0_0_2 = to_unsigned(16#0022#, 16) ELSE
      sbox(34) WHEN out0_0_2 = to_unsigned(16#0023#, 16) ELSE
      sbox(35) WHEN out0_0_2 = to_unsigned(16#0024#, 16) ELSE
      sbox(36) WHEN out0_0_2 = to_unsigned(16#0025#, 16) ELSE
      sbox(37) WHEN out0_0_2 = to_unsigned(16#0026#, 16) ELSE
      sbox(38) WHEN out0_0_2 = to_unsigned(16#0027#, 16) ELSE
      sbox(39) WHEN out0_0_2 = to_unsigned(16#0028#, 16) ELSE
      sbox(40) WHEN out0_0_2 = to_unsigned(16#0029#, 16) ELSE
      sbox(41) WHEN out0_0_2 = to_unsigned(16#002A#, 16) ELSE
      sbox(42) WHEN out0_0_2 = to_unsigned(16#002B#, 16) ELSE
      sbox(43) WHEN out0_0_2 = to_unsigned(16#002C#, 16) ELSE
      sbox(44) WHEN out0_0_2 = to_unsigned(16#002D#, 16) ELSE
      sbox(45) WHEN out0_0_2 = to_unsigned(16#002E#, 16) ELSE
      sbox(46) WHEN out0_0_2 = to_unsigned(16#002F#, 16) ELSE
      sbox(47) WHEN out0_0_2 = to_unsigned(16#0030#, 16) ELSE
      sbox(48) WHEN out0_0_2 = to_unsigned(16#0031#, 16) ELSE
      sbox(49) WHEN out0_0_2 = to_unsigned(16#0032#, 16) ELSE
      sbox(50) WHEN out0_0_2 = to_unsigned(16#0033#, 16) ELSE
      sbox(51) WHEN out0_0_2 = to_unsigned(16#0034#, 16) ELSE
      sbox(52) WHEN out0_0_2 = to_unsigned(16#0035#, 16) ELSE
      sbox(53) WHEN out0_0_2 = to_unsigned(16#0036#, 16) ELSE
      sbox(54) WHEN out0_0_2 = to_unsigned(16#0037#, 16) ELSE
      sbox(55) WHEN out0_0_2 = to_unsigned(16#0038#, 16) ELSE
      sbox(56) WHEN out0_0_2 = to_unsigned(16#0039#, 16) ELSE
      sbox(57) WHEN out0_0_2 = to_unsigned(16#003A#, 16) ELSE
      sbox(58) WHEN out0_0_2 = to_unsigned(16#003B#, 16) ELSE
      sbox(59) WHEN out0_0_2 = to_unsigned(16#003C#, 16) ELSE
      sbox(60) WHEN out0_0_2 = to_unsigned(16#003D#, 16) ELSE
      sbox(61) WHEN out0_0_2 = to_unsigned(16#003E#, 16) ELSE
      sbox(62) WHEN out0_0_2 = to_unsigned(16#003F#, 16) ELSE
      sbox(63) WHEN out0_0_2 = to_unsigned(16#0040#, 16) ELSE
      sbox(64) WHEN out0_0_2 = to_unsigned(16#0041#, 16) ELSE
      sbox(65) WHEN out0_0_2 = to_unsigned(16#0042#, 16) ELSE
      sbox(66) WHEN out0_0_2 = to_unsigned(16#0043#, 16) ELSE
      sbox(67) WHEN out0_0_2 = to_unsigned(16#0044#, 16) ELSE
      sbox(68) WHEN out0_0_2 = to_unsigned(16#0045#, 16) ELSE
      sbox(69) WHEN out0_0_2 = to_unsigned(16#0046#, 16) ELSE
      sbox(70) WHEN out0_0_2 = to_unsigned(16#0047#, 16) ELSE
      sbox(71) WHEN out0_0_2 = to_unsigned(16#0048#, 16) ELSE
      sbox(72) WHEN out0_0_2 = to_unsigned(16#0049#, 16) ELSE
      sbox(73) WHEN out0_0_2 = to_unsigned(16#004A#, 16) ELSE
      sbox(74) WHEN out0_0_2 = to_unsigned(16#004B#, 16) ELSE
      sbox(75) WHEN out0_0_2 = to_unsigned(16#004C#, 16) ELSE
      sbox(76) WHEN out0_0_2 = to_unsigned(16#004D#, 16) ELSE
      sbox(77) WHEN out0_0_2 = to_unsigned(16#004E#, 16) ELSE
      sbox(78) WHEN out0_0_2 = to_unsigned(16#004F#, 16) ELSE
      sbox(79) WHEN out0_0_2 = to_unsigned(16#0050#, 16) ELSE
      sbox(80) WHEN out0_0_2 = to_unsigned(16#0051#, 16) ELSE
      sbox(81) WHEN out0_0_2 = to_unsigned(16#0052#, 16) ELSE
      sbox(82) WHEN out0_0_2 = to_unsigned(16#0053#, 16) ELSE
      sbox(83) WHEN out0_0_2 = to_unsigned(16#0054#, 16) ELSE
      sbox(84) WHEN out0_0_2 = to_unsigned(16#0055#, 16) ELSE
      sbox(85) WHEN out0_0_2 = to_unsigned(16#0056#, 16) ELSE
      sbox(86) WHEN out0_0_2 = to_unsigned(16#0057#, 16) ELSE
      sbox(87) WHEN out0_0_2 = to_unsigned(16#0058#, 16) ELSE
      sbox(88) WHEN out0_0_2 = to_unsigned(16#0059#, 16) ELSE
      sbox(89) WHEN out0_0_2 = to_unsigned(16#005A#, 16) ELSE
      sbox(90) WHEN out0_0_2 = to_unsigned(16#005B#, 16) ELSE
      sbox(91) WHEN out0_0_2 = to_unsigned(16#005C#, 16) ELSE
      sbox(92) WHEN out0_0_2 = to_unsigned(16#005D#, 16) ELSE
      sbox(93) WHEN out0_0_2 = to_unsigned(16#005E#, 16) ELSE
      sbox(94) WHEN out0_0_2 = to_unsigned(16#005F#, 16) ELSE
      sbox(95) WHEN out0_0_2 = to_unsigned(16#0060#, 16) ELSE
      sbox(96) WHEN out0_0_2 = to_unsigned(16#0061#, 16) ELSE
      sbox(97) WHEN out0_0_2 = to_unsigned(16#0062#, 16) ELSE
      sbox(98) WHEN out0_0_2 = to_unsigned(16#0063#, 16) ELSE
      sbox(99) WHEN out0_0_2 = to_unsigned(16#0064#, 16) ELSE
      sbox(100) WHEN out0_0_2 = to_unsigned(16#0065#, 16) ELSE
      sbox(101) WHEN out0_0_2 = to_unsigned(16#0066#, 16) ELSE
      sbox(102) WHEN out0_0_2 = to_unsigned(16#0067#, 16) ELSE
      sbox(103) WHEN out0_0_2 = to_unsigned(16#0068#, 16) ELSE
      sbox(104) WHEN out0_0_2 = to_unsigned(16#0069#, 16) ELSE
      sbox(105) WHEN out0_0_2 = to_unsigned(16#006A#, 16) ELSE
      sbox(106) WHEN out0_0_2 = to_unsigned(16#006B#, 16) ELSE
      sbox(107) WHEN out0_0_2 = to_unsigned(16#006C#, 16) ELSE
      sbox(108) WHEN out0_0_2 = to_unsigned(16#006D#, 16) ELSE
      sbox(109) WHEN out0_0_2 = to_unsigned(16#006E#, 16) ELSE
      sbox(110) WHEN out0_0_2 = to_unsigned(16#006F#, 16) ELSE
      sbox(111) WHEN out0_0_2 = to_unsigned(16#0070#, 16) ELSE
      sbox(112) WHEN out0_0_2 = to_unsigned(16#0071#, 16) ELSE
      sbox(113) WHEN out0_0_2 = to_unsigned(16#0072#, 16) ELSE
      sbox(114) WHEN out0_0_2 = to_unsigned(16#0073#, 16) ELSE
      sbox(115) WHEN out0_0_2 = to_unsigned(16#0074#, 16) ELSE
      sbox(116) WHEN out0_0_2 = to_unsigned(16#0075#, 16) ELSE
      sbox(117) WHEN out0_0_2 = to_unsigned(16#0076#, 16) ELSE
      sbox(118) WHEN out0_0_2 = to_unsigned(16#0077#, 16) ELSE
      sbox(119) WHEN out0_0_2 = to_unsigned(16#0078#, 16) ELSE
      sbox(120) WHEN out0_0_2 = to_unsigned(16#0079#, 16) ELSE
      sbox(121) WHEN out0_0_2 = to_unsigned(16#007A#, 16) ELSE
      sbox(122) WHEN out0_0_2 = to_unsigned(16#007B#, 16) ELSE
      sbox(123) WHEN out0_0_2 = to_unsigned(16#007C#, 16) ELSE
      sbox(124) WHEN out0_0_2 = to_unsigned(16#007D#, 16) ELSE
      sbox(125) WHEN out0_0_2 = to_unsigned(16#007E#, 16) ELSE
      sbox(126) WHEN out0_0_2 = to_unsigned(16#007F#, 16) ELSE
      sbox(127) WHEN out0_0_2 = to_unsigned(16#0080#, 16) ELSE
      sbox(128) WHEN out0_0_2 = to_unsigned(16#0081#, 16) ELSE
      sbox(129) WHEN out0_0_2 = to_unsigned(16#0082#, 16) ELSE
      sbox(130) WHEN out0_0_2 = to_unsigned(16#0083#, 16) ELSE
      sbox(131) WHEN out0_0_2 = to_unsigned(16#0084#, 16) ELSE
      sbox(132) WHEN out0_0_2 = to_unsigned(16#0085#, 16) ELSE
      sbox(133) WHEN out0_0_2 = to_unsigned(16#0086#, 16) ELSE
      sbox(134) WHEN out0_0_2 = to_unsigned(16#0087#, 16) ELSE
      sbox(135) WHEN out0_0_2 = to_unsigned(16#0088#, 16) ELSE
      sbox(136) WHEN out0_0_2 = to_unsigned(16#0089#, 16) ELSE
      sbox(137) WHEN out0_0_2 = to_unsigned(16#008A#, 16) ELSE
      sbox(138) WHEN out0_0_2 = to_unsigned(16#008B#, 16) ELSE
      sbox(139) WHEN out0_0_2 = to_unsigned(16#008C#, 16) ELSE
      sbox(140) WHEN out0_0_2 = to_unsigned(16#008D#, 16) ELSE
      sbox(141) WHEN out0_0_2 = to_unsigned(16#008E#, 16) ELSE
      sbox(142) WHEN out0_0_2 = to_unsigned(16#008F#, 16) ELSE
      sbox(143) WHEN out0_0_2 = to_unsigned(16#0090#, 16) ELSE
      sbox(144) WHEN out0_0_2 = to_unsigned(16#0091#, 16) ELSE
      sbox(145) WHEN out0_0_2 = to_unsigned(16#0092#, 16) ELSE
      sbox(146) WHEN out0_0_2 = to_unsigned(16#0093#, 16) ELSE
      sbox(147) WHEN out0_0_2 = to_unsigned(16#0094#, 16) ELSE
      sbox(148) WHEN out0_0_2 = to_unsigned(16#0095#, 16) ELSE
      sbox(149) WHEN out0_0_2 = to_unsigned(16#0096#, 16) ELSE
      sbox(150) WHEN out0_0_2 = to_unsigned(16#0097#, 16) ELSE
      sbox(151) WHEN out0_0_2 = to_unsigned(16#0098#, 16) ELSE
      sbox(152) WHEN out0_0_2 = to_unsigned(16#0099#, 16) ELSE
      sbox(153) WHEN out0_0_2 = to_unsigned(16#009A#, 16) ELSE
      sbox(154) WHEN out0_0_2 = to_unsigned(16#009B#, 16) ELSE
      sbox(155) WHEN out0_0_2 = to_unsigned(16#009C#, 16) ELSE
      sbox(156) WHEN out0_0_2 = to_unsigned(16#009D#, 16) ELSE
      sbox(157) WHEN out0_0_2 = to_unsigned(16#009E#, 16) ELSE
      sbox(158) WHEN out0_0_2 = to_unsigned(16#009F#, 16) ELSE
      sbox(159) WHEN out0_0_2 = to_unsigned(16#00A0#, 16) ELSE
      sbox(160) WHEN out0_0_2 = to_unsigned(16#00A1#, 16) ELSE
      sbox(161) WHEN out0_0_2 = to_unsigned(16#00A2#, 16) ELSE
      sbox(162) WHEN out0_0_2 = to_unsigned(16#00A3#, 16) ELSE
      sbox(163) WHEN out0_0_2 = to_unsigned(16#00A4#, 16) ELSE
      sbox(164) WHEN out0_0_2 = to_unsigned(16#00A5#, 16) ELSE
      sbox(165) WHEN out0_0_2 = to_unsigned(16#00A6#, 16) ELSE
      sbox(166) WHEN out0_0_2 = to_unsigned(16#00A7#, 16) ELSE
      sbox(167) WHEN out0_0_2 = to_unsigned(16#00A8#, 16) ELSE
      sbox(168) WHEN out0_0_2 = to_unsigned(16#00A9#, 16) ELSE
      sbox(169) WHEN out0_0_2 = to_unsigned(16#00AA#, 16) ELSE
      sbox(170) WHEN out0_0_2 = to_unsigned(16#00AB#, 16) ELSE
      sbox(171) WHEN out0_0_2 = to_unsigned(16#00AC#, 16) ELSE
      sbox(172) WHEN out0_0_2 = to_unsigned(16#00AD#, 16) ELSE
      sbox(173) WHEN out0_0_2 = to_unsigned(16#00AE#, 16) ELSE
      sbox(174) WHEN out0_0_2 = to_unsigned(16#00AF#, 16) ELSE
      sbox(175) WHEN out0_0_2 = to_unsigned(16#00B0#, 16) ELSE
      sbox(176) WHEN out0_0_2 = to_unsigned(16#00B1#, 16) ELSE
      sbox(177) WHEN out0_0_2 = to_unsigned(16#00B2#, 16) ELSE
      sbox(178) WHEN out0_0_2 = to_unsigned(16#00B3#, 16) ELSE
      sbox(179) WHEN out0_0_2 = to_unsigned(16#00B4#, 16) ELSE
      sbox(180) WHEN out0_0_2 = to_unsigned(16#00B5#, 16) ELSE
      sbox(181) WHEN out0_0_2 = to_unsigned(16#00B6#, 16) ELSE
      sbox(182) WHEN out0_0_2 = to_unsigned(16#00B7#, 16) ELSE
      sbox(183) WHEN out0_0_2 = to_unsigned(16#00B8#, 16) ELSE
      sbox(184) WHEN out0_0_2 = to_unsigned(16#00B9#, 16) ELSE
      sbox(185) WHEN out0_0_2 = to_unsigned(16#00BA#, 16) ELSE
      sbox(186) WHEN out0_0_2 = to_unsigned(16#00BB#, 16) ELSE
      sbox(187) WHEN out0_0_2 = to_unsigned(16#00BC#, 16) ELSE
      sbox(188) WHEN out0_0_2 = to_unsigned(16#00BD#, 16) ELSE
      sbox(189) WHEN out0_0_2 = to_unsigned(16#00BE#, 16) ELSE
      sbox(190) WHEN out0_0_2 = to_unsigned(16#00BF#, 16) ELSE
      sbox(191) WHEN out0_0_2 = to_unsigned(16#00C0#, 16) ELSE
      sbox(192) WHEN out0_0_2 = to_unsigned(16#00C1#, 16) ELSE
      sbox(193) WHEN out0_0_2 = to_unsigned(16#00C2#, 16) ELSE
      sbox(194) WHEN out0_0_2 = to_unsigned(16#00C3#, 16) ELSE
      sbox(195) WHEN out0_0_2 = to_unsigned(16#00C4#, 16) ELSE
      sbox(196) WHEN out0_0_2 = to_unsigned(16#00C5#, 16) ELSE
      sbox(197) WHEN out0_0_2 = to_unsigned(16#00C6#, 16) ELSE
      sbox(198) WHEN out0_0_2 = to_unsigned(16#00C7#, 16) ELSE
      sbox(199) WHEN out0_0_2 = to_unsigned(16#00C8#, 16) ELSE
      sbox(200) WHEN out0_0_2 = to_unsigned(16#00C9#, 16) ELSE
      sbox(201) WHEN out0_0_2 = to_unsigned(16#00CA#, 16) ELSE
      sbox(202) WHEN out0_0_2 = to_unsigned(16#00CB#, 16) ELSE
      sbox(203) WHEN out0_0_2 = to_unsigned(16#00CC#, 16) ELSE
      sbox(204) WHEN out0_0_2 = to_unsigned(16#00CD#, 16) ELSE
      sbox(205) WHEN out0_0_2 = to_unsigned(16#00CE#, 16) ELSE
      sbox(206) WHEN out0_0_2 = to_unsigned(16#00CF#, 16) ELSE
      sbox(207) WHEN out0_0_2 = to_unsigned(16#00D0#, 16) ELSE
      sbox(208) WHEN out0_0_2 = to_unsigned(16#00D1#, 16) ELSE
      sbox(209) WHEN out0_0_2 = to_unsigned(16#00D2#, 16) ELSE
      sbox(210) WHEN out0_0_2 = to_unsigned(16#00D3#, 16) ELSE
      sbox(211) WHEN out0_0_2 = to_unsigned(16#00D4#, 16) ELSE
      sbox(212) WHEN out0_0_2 = to_unsigned(16#00D5#, 16) ELSE
      sbox(213) WHEN out0_0_2 = to_unsigned(16#00D6#, 16) ELSE
      sbox(214) WHEN out0_0_2 = to_unsigned(16#00D7#, 16) ELSE
      sbox(215) WHEN out0_0_2 = to_unsigned(16#00D8#, 16) ELSE
      sbox(216) WHEN out0_0_2 = to_unsigned(16#00D9#, 16) ELSE
      sbox(217) WHEN out0_0_2 = to_unsigned(16#00DA#, 16) ELSE
      sbox(218) WHEN out0_0_2 = to_unsigned(16#00DB#, 16) ELSE
      sbox(219) WHEN out0_0_2 = to_unsigned(16#00DC#, 16) ELSE
      sbox(220) WHEN out0_0_2 = to_unsigned(16#00DD#, 16) ELSE
      sbox(221) WHEN out0_0_2 = to_unsigned(16#00DE#, 16) ELSE
      sbox(222) WHEN out0_0_2 = to_unsigned(16#00DF#, 16) ELSE
      sbox(223) WHEN out0_0_2 = to_unsigned(16#00E0#, 16) ELSE
      sbox(224) WHEN out0_0_2 = to_unsigned(16#00E1#, 16) ELSE
      sbox(225) WHEN out0_0_2 = to_unsigned(16#00E2#, 16) ELSE
      sbox(226) WHEN out0_0_2 = to_unsigned(16#00E3#, 16) ELSE
      sbox(227) WHEN out0_0_2 = to_unsigned(16#00E4#, 16) ELSE
      sbox(228) WHEN out0_0_2 = to_unsigned(16#00E5#, 16) ELSE
      sbox(229) WHEN out0_0_2 = to_unsigned(16#00E6#, 16) ELSE
      sbox(230) WHEN out0_0_2 = to_unsigned(16#00E7#, 16) ELSE
      sbox(231) WHEN out0_0_2 = to_unsigned(16#00E8#, 16) ELSE
      sbox(232) WHEN out0_0_2 = to_unsigned(16#00E9#, 16) ELSE
      sbox(233) WHEN out0_0_2 = to_unsigned(16#00EA#, 16) ELSE
      sbox(234) WHEN out0_0_2 = to_unsigned(16#00EB#, 16) ELSE
      sbox(235) WHEN out0_0_2 = to_unsigned(16#00EC#, 16) ELSE
      sbox(236) WHEN out0_0_2 = to_unsigned(16#00ED#, 16) ELSE
      sbox(237) WHEN out0_0_2 = to_unsigned(16#00EE#, 16) ELSE
      sbox(238) WHEN out0_0_2 = to_unsigned(16#00EF#, 16) ELSE
      sbox(239) WHEN out0_0_2 = to_unsigned(16#00F0#, 16) ELSE
      sbox(240) WHEN out0_0_2 = to_unsigned(16#00F1#, 16) ELSE
      sbox(241) WHEN out0_0_2 = to_unsigned(16#00F2#, 16) ELSE
      sbox(242) WHEN out0_0_2 = to_unsigned(16#00F3#, 16) ELSE
      sbox(243) WHEN out0_0_2 = to_unsigned(16#00F4#, 16) ELSE
      sbox(244) WHEN out0_0_2 = to_unsigned(16#00F5#, 16) ELSE
      sbox(245) WHEN out0_0_2 = to_unsigned(16#00F6#, 16) ELSE
      sbox(246) WHEN out0_0_2 = to_unsigned(16#00F7#, 16) ELSE
      sbox(247) WHEN out0_0_2 = to_unsigned(16#00F8#, 16) ELSE
      sbox(248) WHEN out0_0_2 = to_unsigned(16#00F9#, 16) ELSE
      sbox(249) WHEN out0_0_2 = to_unsigned(16#00FA#, 16) ELSE
      sbox(250) WHEN out0_0_2 = to_unsigned(16#00FB#, 16) ELSE
      sbox(251) WHEN out0_0_2 = to_unsigned(16#00FC#, 16) ELSE
      sbox(252) WHEN out0_0_2 = to_unsigned(16#00FD#, 16) ELSE
      sbox(253) WHEN out0_0_2 = to_unsigned(16#00FE#, 16) ELSE
      sbox(254) WHEN out0_0_2 = to_unsigned(16#00FF#, 16) ELSE
      sbox(255);

  s_s_3(0) <= s_0;
  s_s_3(1) <= s_5;
  s_s_3(2) <= s_10;
  s_s_3(3) <= s_15;
  s_s_3(4) <= s_4;
  s_s_3(5) <= s_9;
  s_s_3(6) <= s_14;
  s_s_3(7) <= s_3;
  s_s_3(8) <= s_8;
  s_s_3(9) <= s_13;
  s_s_3(10) <= s_2;
  s_s_3(11) <= s_7;
  s_s_3(12) <= s_12;
  s_s_3(13) <= s_1;
  s_s_3(14) <= s_6;
  s_s_3(15) <= s_11;

  
  out0_127 <= gmul2_15(0) WHEN s_15_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_15(1) WHEN s_15_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_15(2) WHEN s_15_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_15(3) WHEN s_15_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_15(4) WHEN s_15_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_15(5) WHEN s_15_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_15(6) WHEN s_15_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_15(7) WHEN s_15_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_15(8) WHEN s_15_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_15(9) WHEN s_15_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_15(10) WHEN s_15_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_15(11) WHEN s_15_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_15(12) WHEN s_15_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_15(13) WHEN s_15_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_15(14) WHEN s_15_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_15(15) WHEN s_15_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_15(16) WHEN s_15_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_15(17) WHEN s_15_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_15(18) WHEN s_15_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_15(19) WHEN s_15_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_15(20) WHEN s_15_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_15(21) WHEN s_15_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_15(22) WHEN s_15_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_15(23) WHEN s_15_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_15(24) WHEN s_15_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_15(25) WHEN s_15_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_15(26) WHEN s_15_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_15(27) WHEN s_15_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_15(28) WHEN s_15_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_15(29) WHEN s_15_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_15(30) WHEN s_15_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_15(31) WHEN s_15_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_15(32) WHEN s_15_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_15(33) WHEN s_15_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_15(34) WHEN s_15_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_15(35) WHEN s_15_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_15(36) WHEN s_15_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_15(37) WHEN s_15_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_15(38) WHEN s_15_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_15(39) WHEN s_15_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_15(40) WHEN s_15_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_15(41) WHEN s_15_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_15(42) WHEN s_15_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_15(43) WHEN s_15_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_15(44) WHEN s_15_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_15(45) WHEN s_15_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_15(46) WHEN s_15_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_15(47) WHEN s_15_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_15(48) WHEN s_15_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_15(49) WHEN s_15_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_15(50) WHEN s_15_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_15(51) WHEN s_15_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_15(52) WHEN s_15_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_15(53) WHEN s_15_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_15(54) WHEN s_15_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_15(55) WHEN s_15_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_15(56) WHEN s_15_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_15(57) WHEN s_15_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_15(58) WHEN s_15_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_15(59) WHEN s_15_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_15(60) WHEN s_15_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_15(61) WHEN s_15_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_15(62) WHEN s_15_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_15(63) WHEN s_15_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_15(64) WHEN s_15_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_15(65) WHEN s_15_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_15(66) WHEN s_15_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_15(67) WHEN s_15_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_15(68) WHEN s_15_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_15(69) WHEN s_15_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_15(70) WHEN s_15_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_15(71) WHEN s_15_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_15(72) WHEN s_15_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_15(73) WHEN s_15_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_15(74) WHEN s_15_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_15(75) WHEN s_15_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_15(76) WHEN s_15_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_15(77) WHEN s_15_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_15(78) WHEN s_15_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_15(79) WHEN s_15_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_15(80) WHEN s_15_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_15(81) WHEN s_15_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_15(82) WHEN s_15_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_15(83) WHEN s_15_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_15(84) WHEN s_15_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_15(85) WHEN s_15_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_15(86) WHEN s_15_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_15(87) WHEN s_15_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_15(88) WHEN s_15_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_15(89) WHEN s_15_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_15(90) WHEN s_15_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_15(91) WHEN s_15_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_15(92) WHEN s_15_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_15(93) WHEN s_15_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_15(94) WHEN s_15_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_15(95) WHEN s_15_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_15(96) WHEN s_15_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_15(97) WHEN s_15_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_15(98) WHEN s_15_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_15(99) WHEN s_15_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_15(100) WHEN s_15_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_15(101) WHEN s_15_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_15(102) WHEN s_15_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_15(103) WHEN s_15_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_15(104) WHEN s_15_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_15(105) WHEN s_15_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_15(106) WHEN s_15_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_15(107) WHEN s_15_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_15(108) WHEN s_15_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_15(109) WHEN s_15_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_15(110) WHEN s_15_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_15(111) WHEN s_15_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_15(112) WHEN s_15_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_15(113) WHEN s_15_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_15(114) WHEN s_15_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_15(115) WHEN s_15_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_15(116) WHEN s_15_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_15(117) WHEN s_15_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_15(118) WHEN s_15_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_15(119) WHEN s_15_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_15(120) WHEN s_15_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_15(121) WHEN s_15_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_15(122) WHEN s_15_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_15(123) WHEN s_15_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_15(124) WHEN s_15_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_15(125) WHEN s_15_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_15(126) WHEN s_15_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_15(127) WHEN s_15_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_15(128) WHEN s_15_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_15(129) WHEN s_15_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_15(130) WHEN s_15_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_15(131) WHEN s_15_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_15(132) WHEN s_15_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_15(133) WHEN s_15_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_15(134) WHEN s_15_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_15(135) WHEN s_15_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_15(136) WHEN s_15_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_15(137) WHEN s_15_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_15(138) WHEN s_15_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_15(139) WHEN s_15_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_15(140) WHEN s_15_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_15(141) WHEN s_15_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_15(142) WHEN s_15_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_15(143) WHEN s_15_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_15(144) WHEN s_15_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_15(145) WHEN s_15_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_15(146) WHEN s_15_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_15(147) WHEN s_15_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_15(148) WHEN s_15_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_15(149) WHEN s_15_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_15(150) WHEN s_15_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_15(151) WHEN s_15_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_15(152) WHEN s_15_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_15(153) WHEN s_15_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_15(154) WHEN s_15_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_15(155) WHEN s_15_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_15(156) WHEN s_15_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_15(157) WHEN s_15_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_15(158) WHEN s_15_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_15(159) WHEN s_15_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_15(160) WHEN s_15_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_15(161) WHEN s_15_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_15(162) WHEN s_15_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_15(163) WHEN s_15_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_15(164) WHEN s_15_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_15(165) WHEN s_15_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_15(166) WHEN s_15_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_15(167) WHEN s_15_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_15(168) WHEN s_15_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_15(169) WHEN s_15_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_15(170) WHEN s_15_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_15(171) WHEN s_15_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_15(172) WHEN s_15_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_15(173) WHEN s_15_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_15(174) WHEN s_15_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_15(175) WHEN s_15_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_15(176) WHEN s_15_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_15(177) WHEN s_15_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_15(178) WHEN s_15_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_15(179) WHEN s_15_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_15(180) WHEN s_15_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_15(181) WHEN s_15_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_15(182) WHEN s_15_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_15(183) WHEN s_15_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_15(184) WHEN s_15_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_15(185) WHEN s_15_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_15(186) WHEN s_15_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_15(187) WHEN s_15_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_15(188) WHEN s_15_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_15(189) WHEN s_15_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_15(190) WHEN s_15_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_15(191) WHEN s_15_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_15(192) WHEN s_15_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_15(193) WHEN s_15_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_15(194) WHEN s_15_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_15(195) WHEN s_15_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_15(196) WHEN s_15_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_15(197) WHEN s_15_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_15(198) WHEN s_15_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_15(199) WHEN s_15_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_15(200) WHEN s_15_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_15(201) WHEN s_15_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_15(202) WHEN s_15_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_15(203) WHEN s_15_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_15(204) WHEN s_15_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_15(205) WHEN s_15_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_15(206) WHEN s_15_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_15(207) WHEN s_15_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_15(208) WHEN s_15_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_15(209) WHEN s_15_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_15(210) WHEN s_15_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_15(211) WHEN s_15_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_15(212) WHEN s_15_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_15(213) WHEN s_15_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_15(214) WHEN s_15_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_15(215) WHEN s_15_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_15(216) WHEN s_15_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_15(217) WHEN s_15_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_15(218) WHEN s_15_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_15(219) WHEN s_15_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_15(220) WHEN s_15_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_15(221) WHEN s_15_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_15(222) WHEN s_15_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_15(223) WHEN s_15_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_15(224) WHEN s_15_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_15(225) WHEN s_15_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_15(226) WHEN s_15_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_15(227) WHEN s_15_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_15(228) WHEN s_15_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_15(229) WHEN s_15_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_15(230) WHEN s_15_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_15(231) WHEN s_15_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_15(232) WHEN s_15_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_15(233) WHEN s_15_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_15(234) WHEN s_15_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_15(235) WHEN s_15_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_15(236) WHEN s_15_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_15(237) WHEN s_15_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_15(238) WHEN s_15_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_15(239) WHEN s_15_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_15(240) WHEN s_15_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_15(241) WHEN s_15_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_15(242) WHEN s_15_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_15(243) WHEN s_15_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_15(244) WHEN s_15_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_15(245) WHEN s_15_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_15(246) WHEN s_15_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_15(247) WHEN s_15_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_15(248) WHEN s_15_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_15(249) WHEN s_15_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_15(250) WHEN s_15_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_15(251) WHEN s_15_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_15(252) WHEN s_15_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_15(253) WHEN s_15_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_15(254) WHEN s_15_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_15(255);

  
  out0_128 <= gmul3_15(0) WHEN s_12_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_15(1) WHEN s_12_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_15(2) WHEN s_12_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_15(3) WHEN s_12_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_15(4) WHEN s_12_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_15(5) WHEN s_12_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_15(6) WHEN s_12_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_15(7) WHEN s_12_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_15(8) WHEN s_12_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_15(9) WHEN s_12_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_15(10) WHEN s_12_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_15(11) WHEN s_12_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_15(12) WHEN s_12_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_15(13) WHEN s_12_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_15(14) WHEN s_12_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_15(15) WHEN s_12_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_15(16) WHEN s_12_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_15(17) WHEN s_12_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_15(18) WHEN s_12_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_15(19) WHEN s_12_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_15(20) WHEN s_12_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_15(21) WHEN s_12_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_15(22) WHEN s_12_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_15(23) WHEN s_12_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_15(24) WHEN s_12_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_15(25) WHEN s_12_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_15(26) WHEN s_12_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_15(27) WHEN s_12_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_15(28) WHEN s_12_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_15(29) WHEN s_12_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_15(30) WHEN s_12_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_15(31) WHEN s_12_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_15(32) WHEN s_12_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_15(33) WHEN s_12_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_15(34) WHEN s_12_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_15(35) WHEN s_12_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_15(36) WHEN s_12_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_15(37) WHEN s_12_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_15(38) WHEN s_12_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_15(39) WHEN s_12_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_15(40) WHEN s_12_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_15(41) WHEN s_12_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_15(42) WHEN s_12_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_15(43) WHEN s_12_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_15(44) WHEN s_12_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_15(45) WHEN s_12_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_15(46) WHEN s_12_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_15(47) WHEN s_12_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_15(48) WHEN s_12_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_15(49) WHEN s_12_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_15(50) WHEN s_12_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_15(51) WHEN s_12_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_15(52) WHEN s_12_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_15(53) WHEN s_12_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_15(54) WHEN s_12_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_15(55) WHEN s_12_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_15(56) WHEN s_12_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_15(57) WHEN s_12_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_15(58) WHEN s_12_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_15(59) WHEN s_12_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_15(60) WHEN s_12_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_15(61) WHEN s_12_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_15(62) WHEN s_12_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_15(63) WHEN s_12_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_15(64) WHEN s_12_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_15(65) WHEN s_12_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_15(66) WHEN s_12_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_15(67) WHEN s_12_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_15(68) WHEN s_12_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_15(69) WHEN s_12_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_15(70) WHEN s_12_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_15(71) WHEN s_12_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_15(72) WHEN s_12_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_15(73) WHEN s_12_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_15(74) WHEN s_12_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_15(75) WHEN s_12_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_15(76) WHEN s_12_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_15(77) WHEN s_12_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_15(78) WHEN s_12_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_15(79) WHEN s_12_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_15(80) WHEN s_12_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_15(81) WHEN s_12_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_15(82) WHEN s_12_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_15(83) WHEN s_12_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_15(84) WHEN s_12_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_15(85) WHEN s_12_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_15(86) WHEN s_12_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_15(87) WHEN s_12_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_15(88) WHEN s_12_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_15(89) WHEN s_12_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_15(90) WHEN s_12_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_15(91) WHEN s_12_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_15(92) WHEN s_12_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_15(93) WHEN s_12_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_15(94) WHEN s_12_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_15(95) WHEN s_12_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_15(96) WHEN s_12_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_15(97) WHEN s_12_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_15(98) WHEN s_12_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_15(99) WHEN s_12_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_15(100) WHEN s_12_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_15(101) WHEN s_12_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_15(102) WHEN s_12_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_15(103) WHEN s_12_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_15(104) WHEN s_12_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_15(105) WHEN s_12_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_15(106) WHEN s_12_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_15(107) WHEN s_12_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_15(108) WHEN s_12_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_15(109) WHEN s_12_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_15(110) WHEN s_12_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_15(111) WHEN s_12_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_15(112) WHEN s_12_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_15(113) WHEN s_12_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_15(114) WHEN s_12_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_15(115) WHEN s_12_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_15(116) WHEN s_12_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_15(117) WHEN s_12_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_15(118) WHEN s_12_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_15(119) WHEN s_12_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_15(120) WHEN s_12_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_15(121) WHEN s_12_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_15(122) WHEN s_12_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_15(123) WHEN s_12_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_15(124) WHEN s_12_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_15(125) WHEN s_12_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_15(126) WHEN s_12_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_15(127) WHEN s_12_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_15(128) WHEN s_12_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_15(129) WHEN s_12_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_15(130) WHEN s_12_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_15(131) WHEN s_12_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_15(132) WHEN s_12_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_15(133) WHEN s_12_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_15(134) WHEN s_12_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_15(135) WHEN s_12_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_15(136) WHEN s_12_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_15(137) WHEN s_12_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_15(138) WHEN s_12_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_15(139) WHEN s_12_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_15(140) WHEN s_12_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_15(141) WHEN s_12_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_15(142) WHEN s_12_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_15(143) WHEN s_12_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_15(144) WHEN s_12_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_15(145) WHEN s_12_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_15(146) WHEN s_12_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_15(147) WHEN s_12_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_15(148) WHEN s_12_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_15(149) WHEN s_12_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_15(150) WHEN s_12_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_15(151) WHEN s_12_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_15(152) WHEN s_12_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_15(153) WHEN s_12_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_15(154) WHEN s_12_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_15(155) WHEN s_12_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_15(156) WHEN s_12_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_15(157) WHEN s_12_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_15(158) WHEN s_12_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_15(159) WHEN s_12_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_15(160) WHEN s_12_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_15(161) WHEN s_12_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_15(162) WHEN s_12_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_15(163) WHEN s_12_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_15(164) WHEN s_12_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_15(165) WHEN s_12_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_15(166) WHEN s_12_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_15(167) WHEN s_12_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_15(168) WHEN s_12_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_15(169) WHEN s_12_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_15(170) WHEN s_12_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_15(171) WHEN s_12_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_15(172) WHEN s_12_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_15(173) WHEN s_12_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_15(174) WHEN s_12_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_15(175) WHEN s_12_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_15(176) WHEN s_12_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_15(177) WHEN s_12_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_15(178) WHEN s_12_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_15(179) WHEN s_12_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_15(180) WHEN s_12_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_15(181) WHEN s_12_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_15(182) WHEN s_12_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_15(183) WHEN s_12_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_15(184) WHEN s_12_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_15(185) WHEN s_12_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_15(186) WHEN s_12_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_15(187) WHEN s_12_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_15(188) WHEN s_12_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_15(189) WHEN s_12_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_15(190) WHEN s_12_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_15(191) WHEN s_12_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_15(192) WHEN s_12_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_15(193) WHEN s_12_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_15(194) WHEN s_12_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_15(195) WHEN s_12_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_15(196) WHEN s_12_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_15(197) WHEN s_12_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_15(198) WHEN s_12_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_15(199) WHEN s_12_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_15(200) WHEN s_12_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_15(201) WHEN s_12_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_15(202) WHEN s_12_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_15(203) WHEN s_12_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_15(204) WHEN s_12_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_15(205) WHEN s_12_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_15(206) WHEN s_12_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_15(207) WHEN s_12_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_15(208) WHEN s_12_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_15(209) WHEN s_12_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_15(210) WHEN s_12_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_15(211) WHEN s_12_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_15(212) WHEN s_12_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_15(213) WHEN s_12_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_15(214) WHEN s_12_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_15(215) WHEN s_12_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_15(216) WHEN s_12_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_15(217) WHEN s_12_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_15(218) WHEN s_12_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_15(219) WHEN s_12_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_15(220) WHEN s_12_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_15(221) WHEN s_12_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_15(222) WHEN s_12_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_15(223) WHEN s_12_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_15(224) WHEN s_12_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_15(225) WHEN s_12_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_15(226) WHEN s_12_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_15(227) WHEN s_12_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_15(228) WHEN s_12_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_15(229) WHEN s_12_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_15(230) WHEN s_12_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_15(231) WHEN s_12_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_15(232) WHEN s_12_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_15(233) WHEN s_12_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_15(234) WHEN s_12_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_15(235) WHEN s_12_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_15(236) WHEN s_12_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_15(237) WHEN s_12_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_15(238) WHEN s_12_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_15(239) WHEN s_12_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_15(240) WHEN s_12_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_15(241) WHEN s_12_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_15(242) WHEN s_12_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_15(243) WHEN s_12_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_15(244) WHEN s_12_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_15(245) WHEN s_12_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_15(246) WHEN s_12_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_15(247) WHEN s_12_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_15(248) WHEN s_12_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_15(249) WHEN s_12_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_15(250) WHEN s_12_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_15(251) WHEN s_12_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_15(252) WHEN s_12_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_15(253) WHEN s_12_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_15(254) WHEN s_12_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_15(255);

  out0_129 <= out0_128 XOR s_13_1;

  b4 <= out0_129 XOR s_14_1;

  out0_130 <= b4 XOR out0_127;

  
  out0_131 <= gmul3_14(0) WHEN s_15_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_14(1) WHEN s_15_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_14(2) WHEN s_15_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_14(3) WHEN s_15_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_14(4) WHEN s_15_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_14(5) WHEN s_15_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_14(6) WHEN s_15_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_14(7) WHEN s_15_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_14(8) WHEN s_15_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_14(9) WHEN s_15_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_14(10) WHEN s_15_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_14(11) WHEN s_15_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_14(12) WHEN s_15_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_14(13) WHEN s_15_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_14(14) WHEN s_15_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_14(15) WHEN s_15_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_14(16) WHEN s_15_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_14(17) WHEN s_15_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_14(18) WHEN s_15_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_14(19) WHEN s_15_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_14(20) WHEN s_15_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_14(21) WHEN s_15_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_14(22) WHEN s_15_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_14(23) WHEN s_15_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_14(24) WHEN s_15_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_14(25) WHEN s_15_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_14(26) WHEN s_15_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_14(27) WHEN s_15_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_14(28) WHEN s_15_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_14(29) WHEN s_15_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_14(30) WHEN s_15_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_14(31) WHEN s_15_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_14(32) WHEN s_15_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_14(33) WHEN s_15_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_14(34) WHEN s_15_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_14(35) WHEN s_15_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_14(36) WHEN s_15_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_14(37) WHEN s_15_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_14(38) WHEN s_15_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_14(39) WHEN s_15_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_14(40) WHEN s_15_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_14(41) WHEN s_15_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_14(42) WHEN s_15_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_14(43) WHEN s_15_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_14(44) WHEN s_15_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_14(45) WHEN s_15_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_14(46) WHEN s_15_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_14(47) WHEN s_15_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_14(48) WHEN s_15_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_14(49) WHEN s_15_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_14(50) WHEN s_15_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_14(51) WHEN s_15_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_14(52) WHEN s_15_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_14(53) WHEN s_15_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_14(54) WHEN s_15_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_14(55) WHEN s_15_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_14(56) WHEN s_15_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_14(57) WHEN s_15_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_14(58) WHEN s_15_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_14(59) WHEN s_15_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_14(60) WHEN s_15_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_14(61) WHEN s_15_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_14(62) WHEN s_15_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_14(63) WHEN s_15_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_14(64) WHEN s_15_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_14(65) WHEN s_15_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_14(66) WHEN s_15_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_14(67) WHEN s_15_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_14(68) WHEN s_15_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_14(69) WHEN s_15_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_14(70) WHEN s_15_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_14(71) WHEN s_15_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_14(72) WHEN s_15_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_14(73) WHEN s_15_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_14(74) WHEN s_15_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_14(75) WHEN s_15_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_14(76) WHEN s_15_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_14(77) WHEN s_15_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_14(78) WHEN s_15_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_14(79) WHEN s_15_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_14(80) WHEN s_15_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_14(81) WHEN s_15_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_14(82) WHEN s_15_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_14(83) WHEN s_15_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_14(84) WHEN s_15_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_14(85) WHEN s_15_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_14(86) WHEN s_15_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_14(87) WHEN s_15_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_14(88) WHEN s_15_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_14(89) WHEN s_15_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_14(90) WHEN s_15_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_14(91) WHEN s_15_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_14(92) WHEN s_15_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_14(93) WHEN s_15_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_14(94) WHEN s_15_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_14(95) WHEN s_15_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_14(96) WHEN s_15_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_14(97) WHEN s_15_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_14(98) WHEN s_15_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_14(99) WHEN s_15_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_14(100) WHEN s_15_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_14(101) WHEN s_15_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_14(102) WHEN s_15_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_14(103) WHEN s_15_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_14(104) WHEN s_15_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_14(105) WHEN s_15_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_14(106) WHEN s_15_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_14(107) WHEN s_15_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_14(108) WHEN s_15_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_14(109) WHEN s_15_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_14(110) WHEN s_15_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_14(111) WHEN s_15_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_14(112) WHEN s_15_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_14(113) WHEN s_15_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_14(114) WHEN s_15_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_14(115) WHEN s_15_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_14(116) WHEN s_15_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_14(117) WHEN s_15_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_14(118) WHEN s_15_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_14(119) WHEN s_15_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_14(120) WHEN s_15_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_14(121) WHEN s_15_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_14(122) WHEN s_15_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_14(123) WHEN s_15_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_14(124) WHEN s_15_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_14(125) WHEN s_15_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_14(126) WHEN s_15_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_14(127) WHEN s_15_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_14(128) WHEN s_15_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_14(129) WHEN s_15_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_14(130) WHEN s_15_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_14(131) WHEN s_15_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_14(132) WHEN s_15_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_14(133) WHEN s_15_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_14(134) WHEN s_15_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_14(135) WHEN s_15_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_14(136) WHEN s_15_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_14(137) WHEN s_15_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_14(138) WHEN s_15_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_14(139) WHEN s_15_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_14(140) WHEN s_15_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_14(141) WHEN s_15_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_14(142) WHEN s_15_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_14(143) WHEN s_15_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_14(144) WHEN s_15_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_14(145) WHEN s_15_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_14(146) WHEN s_15_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_14(147) WHEN s_15_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_14(148) WHEN s_15_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_14(149) WHEN s_15_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_14(150) WHEN s_15_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_14(151) WHEN s_15_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_14(152) WHEN s_15_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_14(153) WHEN s_15_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_14(154) WHEN s_15_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_14(155) WHEN s_15_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_14(156) WHEN s_15_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_14(157) WHEN s_15_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_14(158) WHEN s_15_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_14(159) WHEN s_15_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_14(160) WHEN s_15_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_14(161) WHEN s_15_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_14(162) WHEN s_15_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_14(163) WHEN s_15_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_14(164) WHEN s_15_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_14(165) WHEN s_15_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_14(166) WHEN s_15_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_14(167) WHEN s_15_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_14(168) WHEN s_15_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_14(169) WHEN s_15_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_14(170) WHEN s_15_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_14(171) WHEN s_15_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_14(172) WHEN s_15_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_14(173) WHEN s_15_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_14(174) WHEN s_15_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_14(175) WHEN s_15_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_14(176) WHEN s_15_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_14(177) WHEN s_15_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_14(178) WHEN s_15_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_14(179) WHEN s_15_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_14(180) WHEN s_15_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_14(181) WHEN s_15_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_14(182) WHEN s_15_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_14(183) WHEN s_15_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_14(184) WHEN s_15_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_14(185) WHEN s_15_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_14(186) WHEN s_15_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_14(187) WHEN s_15_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_14(188) WHEN s_15_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_14(189) WHEN s_15_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_14(190) WHEN s_15_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_14(191) WHEN s_15_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_14(192) WHEN s_15_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_14(193) WHEN s_15_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_14(194) WHEN s_15_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_14(195) WHEN s_15_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_14(196) WHEN s_15_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_14(197) WHEN s_15_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_14(198) WHEN s_15_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_14(199) WHEN s_15_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_14(200) WHEN s_15_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_14(201) WHEN s_15_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_14(202) WHEN s_15_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_14(203) WHEN s_15_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_14(204) WHEN s_15_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_14(205) WHEN s_15_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_14(206) WHEN s_15_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_14(207) WHEN s_15_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_14(208) WHEN s_15_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_14(209) WHEN s_15_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_14(210) WHEN s_15_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_14(211) WHEN s_15_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_14(212) WHEN s_15_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_14(213) WHEN s_15_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_14(214) WHEN s_15_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_14(215) WHEN s_15_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_14(216) WHEN s_15_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_14(217) WHEN s_15_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_14(218) WHEN s_15_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_14(219) WHEN s_15_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_14(220) WHEN s_15_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_14(221) WHEN s_15_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_14(222) WHEN s_15_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_14(223) WHEN s_15_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_14(224) WHEN s_15_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_14(225) WHEN s_15_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_14(226) WHEN s_15_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_14(227) WHEN s_15_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_14(228) WHEN s_15_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_14(229) WHEN s_15_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_14(230) WHEN s_15_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_14(231) WHEN s_15_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_14(232) WHEN s_15_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_14(233) WHEN s_15_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_14(234) WHEN s_15_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_14(235) WHEN s_15_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_14(236) WHEN s_15_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_14(237) WHEN s_15_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_14(238) WHEN s_15_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_14(239) WHEN s_15_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_14(240) WHEN s_15_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_14(241) WHEN s_15_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_14(242) WHEN s_15_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_14(243) WHEN s_15_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_14(244) WHEN s_15_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_14(245) WHEN s_15_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_14(246) WHEN s_15_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_14(247) WHEN s_15_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_14(248) WHEN s_15_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_14(249) WHEN s_15_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_14(250) WHEN s_15_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_14(251) WHEN s_15_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_14(252) WHEN s_15_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_14(253) WHEN s_15_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_14(254) WHEN s_15_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_14(255);

  
  out0_132 <= gmul2_14(0) WHEN s_14_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_14(1) WHEN s_14_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_14(2) WHEN s_14_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_14(3) WHEN s_14_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_14(4) WHEN s_14_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_14(5) WHEN s_14_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_14(6) WHEN s_14_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_14(7) WHEN s_14_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_14(8) WHEN s_14_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_14(9) WHEN s_14_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_14(10) WHEN s_14_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_14(11) WHEN s_14_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_14(12) WHEN s_14_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_14(13) WHEN s_14_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_14(14) WHEN s_14_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_14(15) WHEN s_14_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_14(16) WHEN s_14_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_14(17) WHEN s_14_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_14(18) WHEN s_14_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_14(19) WHEN s_14_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_14(20) WHEN s_14_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_14(21) WHEN s_14_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_14(22) WHEN s_14_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_14(23) WHEN s_14_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_14(24) WHEN s_14_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_14(25) WHEN s_14_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_14(26) WHEN s_14_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_14(27) WHEN s_14_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_14(28) WHEN s_14_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_14(29) WHEN s_14_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_14(30) WHEN s_14_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_14(31) WHEN s_14_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_14(32) WHEN s_14_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_14(33) WHEN s_14_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_14(34) WHEN s_14_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_14(35) WHEN s_14_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_14(36) WHEN s_14_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_14(37) WHEN s_14_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_14(38) WHEN s_14_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_14(39) WHEN s_14_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_14(40) WHEN s_14_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_14(41) WHEN s_14_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_14(42) WHEN s_14_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_14(43) WHEN s_14_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_14(44) WHEN s_14_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_14(45) WHEN s_14_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_14(46) WHEN s_14_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_14(47) WHEN s_14_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_14(48) WHEN s_14_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_14(49) WHEN s_14_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_14(50) WHEN s_14_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_14(51) WHEN s_14_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_14(52) WHEN s_14_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_14(53) WHEN s_14_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_14(54) WHEN s_14_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_14(55) WHEN s_14_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_14(56) WHEN s_14_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_14(57) WHEN s_14_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_14(58) WHEN s_14_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_14(59) WHEN s_14_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_14(60) WHEN s_14_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_14(61) WHEN s_14_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_14(62) WHEN s_14_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_14(63) WHEN s_14_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_14(64) WHEN s_14_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_14(65) WHEN s_14_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_14(66) WHEN s_14_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_14(67) WHEN s_14_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_14(68) WHEN s_14_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_14(69) WHEN s_14_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_14(70) WHEN s_14_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_14(71) WHEN s_14_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_14(72) WHEN s_14_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_14(73) WHEN s_14_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_14(74) WHEN s_14_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_14(75) WHEN s_14_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_14(76) WHEN s_14_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_14(77) WHEN s_14_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_14(78) WHEN s_14_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_14(79) WHEN s_14_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_14(80) WHEN s_14_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_14(81) WHEN s_14_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_14(82) WHEN s_14_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_14(83) WHEN s_14_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_14(84) WHEN s_14_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_14(85) WHEN s_14_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_14(86) WHEN s_14_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_14(87) WHEN s_14_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_14(88) WHEN s_14_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_14(89) WHEN s_14_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_14(90) WHEN s_14_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_14(91) WHEN s_14_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_14(92) WHEN s_14_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_14(93) WHEN s_14_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_14(94) WHEN s_14_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_14(95) WHEN s_14_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_14(96) WHEN s_14_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_14(97) WHEN s_14_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_14(98) WHEN s_14_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_14(99) WHEN s_14_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_14(100) WHEN s_14_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_14(101) WHEN s_14_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_14(102) WHEN s_14_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_14(103) WHEN s_14_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_14(104) WHEN s_14_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_14(105) WHEN s_14_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_14(106) WHEN s_14_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_14(107) WHEN s_14_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_14(108) WHEN s_14_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_14(109) WHEN s_14_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_14(110) WHEN s_14_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_14(111) WHEN s_14_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_14(112) WHEN s_14_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_14(113) WHEN s_14_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_14(114) WHEN s_14_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_14(115) WHEN s_14_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_14(116) WHEN s_14_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_14(117) WHEN s_14_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_14(118) WHEN s_14_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_14(119) WHEN s_14_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_14(120) WHEN s_14_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_14(121) WHEN s_14_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_14(122) WHEN s_14_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_14(123) WHEN s_14_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_14(124) WHEN s_14_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_14(125) WHEN s_14_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_14(126) WHEN s_14_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_14(127) WHEN s_14_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_14(128) WHEN s_14_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_14(129) WHEN s_14_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_14(130) WHEN s_14_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_14(131) WHEN s_14_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_14(132) WHEN s_14_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_14(133) WHEN s_14_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_14(134) WHEN s_14_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_14(135) WHEN s_14_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_14(136) WHEN s_14_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_14(137) WHEN s_14_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_14(138) WHEN s_14_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_14(139) WHEN s_14_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_14(140) WHEN s_14_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_14(141) WHEN s_14_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_14(142) WHEN s_14_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_14(143) WHEN s_14_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_14(144) WHEN s_14_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_14(145) WHEN s_14_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_14(146) WHEN s_14_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_14(147) WHEN s_14_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_14(148) WHEN s_14_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_14(149) WHEN s_14_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_14(150) WHEN s_14_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_14(151) WHEN s_14_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_14(152) WHEN s_14_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_14(153) WHEN s_14_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_14(154) WHEN s_14_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_14(155) WHEN s_14_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_14(156) WHEN s_14_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_14(157) WHEN s_14_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_14(158) WHEN s_14_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_14(159) WHEN s_14_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_14(160) WHEN s_14_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_14(161) WHEN s_14_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_14(162) WHEN s_14_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_14(163) WHEN s_14_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_14(164) WHEN s_14_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_14(165) WHEN s_14_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_14(166) WHEN s_14_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_14(167) WHEN s_14_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_14(168) WHEN s_14_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_14(169) WHEN s_14_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_14(170) WHEN s_14_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_14(171) WHEN s_14_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_14(172) WHEN s_14_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_14(173) WHEN s_14_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_14(174) WHEN s_14_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_14(175) WHEN s_14_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_14(176) WHEN s_14_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_14(177) WHEN s_14_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_14(178) WHEN s_14_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_14(179) WHEN s_14_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_14(180) WHEN s_14_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_14(181) WHEN s_14_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_14(182) WHEN s_14_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_14(183) WHEN s_14_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_14(184) WHEN s_14_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_14(185) WHEN s_14_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_14(186) WHEN s_14_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_14(187) WHEN s_14_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_14(188) WHEN s_14_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_14(189) WHEN s_14_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_14(190) WHEN s_14_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_14(191) WHEN s_14_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_14(192) WHEN s_14_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_14(193) WHEN s_14_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_14(194) WHEN s_14_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_14(195) WHEN s_14_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_14(196) WHEN s_14_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_14(197) WHEN s_14_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_14(198) WHEN s_14_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_14(199) WHEN s_14_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_14(200) WHEN s_14_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_14(201) WHEN s_14_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_14(202) WHEN s_14_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_14(203) WHEN s_14_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_14(204) WHEN s_14_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_14(205) WHEN s_14_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_14(206) WHEN s_14_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_14(207) WHEN s_14_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_14(208) WHEN s_14_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_14(209) WHEN s_14_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_14(210) WHEN s_14_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_14(211) WHEN s_14_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_14(212) WHEN s_14_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_14(213) WHEN s_14_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_14(214) WHEN s_14_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_14(215) WHEN s_14_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_14(216) WHEN s_14_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_14(217) WHEN s_14_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_14(218) WHEN s_14_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_14(219) WHEN s_14_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_14(220) WHEN s_14_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_14(221) WHEN s_14_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_14(222) WHEN s_14_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_14(223) WHEN s_14_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_14(224) WHEN s_14_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_14(225) WHEN s_14_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_14(226) WHEN s_14_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_14(227) WHEN s_14_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_14(228) WHEN s_14_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_14(229) WHEN s_14_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_14(230) WHEN s_14_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_14(231) WHEN s_14_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_14(232) WHEN s_14_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_14(233) WHEN s_14_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_14(234) WHEN s_14_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_14(235) WHEN s_14_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_14(236) WHEN s_14_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_14(237) WHEN s_14_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_14(238) WHEN s_14_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_14(239) WHEN s_14_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_14(240) WHEN s_14_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_14(241) WHEN s_14_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_14(242) WHEN s_14_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_14(243) WHEN s_14_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_14(244) WHEN s_14_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_14(245) WHEN s_14_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_14(246) WHEN s_14_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_14(247) WHEN s_14_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_14(248) WHEN s_14_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_14(249) WHEN s_14_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_14(250) WHEN s_14_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_14(251) WHEN s_14_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_14(252) WHEN s_14_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_14(253) WHEN s_14_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_14(254) WHEN s_14_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_14(255);

  out0_133 <= s_12_1 XOR s_13_1;

  b3 <= out0_133 XOR out0_132;

  out0_134 <= b3 XOR out0_131;

  
  out0_135 <= gmul3_13(0) WHEN s_14_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_13(1) WHEN s_14_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_13(2) WHEN s_14_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_13(3) WHEN s_14_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_13(4) WHEN s_14_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_13(5) WHEN s_14_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_13(6) WHEN s_14_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_13(7) WHEN s_14_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_13(8) WHEN s_14_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_13(9) WHEN s_14_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_13(10) WHEN s_14_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_13(11) WHEN s_14_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_13(12) WHEN s_14_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_13(13) WHEN s_14_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_13(14) WHEN s_14_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_13(15) WHEN s_14_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_13(16) WHEN s_14_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_13(17) WHEN s_14_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_13(18) WHEN s_14_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_13(19) WHEN s_14_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_13(20) WHEN s_14_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_13(21) WHEN s_14_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_13(22) WHEN s_14_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_13(23) WHEN s_14_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_13(24) WHEN s_14_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_13(25) WHEN s_14_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_13(26) WHEN s_14_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_13(27) WHEN s_14_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_13(28) WHEN s_14_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_13(29) WHEN s_14_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_13(30) WHEN s_14_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_13(31) WHEN s_14_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_13(32) WHEN s_14_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_13(33) WHEN s_14_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_13(34) WHEN s_14_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_13(35) WHEN s_14_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_13(36) WHEN s_14_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_13(37) WHEN s_14_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_13(38) WHEN s_14_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_13(39) WHEN s_14_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_13(40) WHEN s_14_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_13(41) WHEN s_14_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_13(42) WHEN s_14_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_13(43) WHEN s_14_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_13(44) WHEN s_14_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_13(45) WHEN s_14_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_13(46) WHEN s_14_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_13(47) WHEN s_14_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_13(48) WHEN s_14_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_13(49) WHEN s_14_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_13(50) WHEN s_14_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_13(51) WHEN s_14_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_13(52) WHEN s_14_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_13(53) WHEN s_14_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_13(54) WHEN s_14_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_13(55) WHEN s_14_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_13(56) WHEN s_14_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_13(57) WHEN s_14_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_13(58) WHEN s_14_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_13(59) WHEN s_14_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_13(60) WHEN s_14_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_13(61) WHEN s_14_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_13(62) WHEN s_14_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_13(63) WHEN s_14_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_13(64) WHEN s_14_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_13(65) WHEN s_14_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_13(66) WHEN s_14_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_13(67) WHEN s_14_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_13(68) WHEN s_14_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_13(69) WHEN s_14_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_13(70) WHEN s_14_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_13(71) WHEN s_14_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_13(72) WHEN s_14_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_13(73) WHEN s_14_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_13(74) WHEN s_14_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_13(75) WHEN s_14_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_13(76) WHEN s_14_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_13(77) WHEN s_14_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_13(78) WHEN s_14_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_13(79) WHEN s_14_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_13(80) WHEN s_14_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_13(81) WHEN s_14_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_13(82) WHEN s_14_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_13(83) WHEN s_14_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_13(84) WHEN s_14_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_13(85) WHEN s_14_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_13(86) WHEN s_14_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_13(87) WHEN s_14_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_13(88) WHEN s_14_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_13(89) WHEN s_14_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_13(90) WHEN s_14_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_13(91) WHEN s_14_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_13(92) WHEN s_14_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_13(93) WHEN s_14_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_13(94) WHEN s_14_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_13(95) WHEN s_14_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_13(96) WHEN s_14_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_13(97) WHEN s_14_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_13(98) WHEN s_14_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_13(99) WHEN s_14_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_13(100) WHEN s_14_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_13(101) WHEN s_14_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_13(102) WHEN s_14_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_13(103) WHEN s_14_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_13(104) WHEN s_14_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_13(105) WHEN s_14_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_13(106) WHEN s_14_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_13(107) WHEN s_14_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_13(108) WHEN s_14_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_13(109) WHEN s_14_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_13(110) WHEN s_14_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_13(111) WHEN s_14_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_13(112) WHEN s_14_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_13(113) WHEN s_14_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_13(114) WHEN s_14_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_13(115) WHEN s_14_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_13(116) WHEN s_14_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_13(117) WHEN s_14_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_13(118) WHEN s_14_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_13(119) WHEN s_14_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_13(120) WHEN s_14_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_13(121) WHEN s_14_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_13(122) WHEN s_14_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_13(123) WHEN s_14_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_13(124) WHEN s_14_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_13(125) WHEN s_14_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_13(126) WHEN s_14_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_13(127) WHEN s_14_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_13(128) WHEN s_14_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_13(129) WHEN s_14_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_13(130) WHEN s_14_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_13(131) WHEN s_14_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_13(132) WHEN s_14_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_13(133) WHEN s_14_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_13(134) WHEN s_14_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_13(135) WHEN s_14_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_13(136) WHEN s_14_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_13(137) WHEN s_14_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_13(138) WHEN s_14_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_13(139) WHEN s_14_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_13(140) WHEN s_14_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_13(141) WHEN s_14_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_13(142) WHEN s_14_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_13(143) WHEN s_14_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_13(144) WHEN s_14_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_13(145) WHEN s_14_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_13(146) WHEN s_14_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_13(147) WHEN s_14_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_13(148) WHEN s_14_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_13(149) WHEN s_14_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_13(150) WHEN s_14_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_13(151) WHEN s_14_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_13(152) WHEN s_14_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_13(153) WHEN s_14_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_13(154) WHEN s_14_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_13(155) WHEN s_14_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_13(156) WHEN s_14_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_13(157) WHEN s_14_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_13(158) WHEN s_14_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_13(159) WHEN s_14_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_13(160) WHEN s_14_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_13(161) WHEN s_14_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_13(162) WHEN s_14_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_13(163) WHEN s_14_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_13(164) WHEN s_14_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_13(165) WHEN s_14_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_13(166) WHEN s_14_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_13(167) WHEN s_14_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_13(168) WHEN s_14_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_13(169) WHEN s_14_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_13(170) WHEN s_14_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_13(171) WHEN s_14_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_13(172) WHEN s_14_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_13(173) WHEN s_14_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_13(174) WHEN s_14_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_13(175) WHEN s_14_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_13(176) WHEN s_14_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_13(177) WHEN s_14_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_13(178) WHEN s_14_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_13(179) WHEN s_14_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_13(180) WHEN s_14_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_13(181) WHEN s_14_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_13(182) WHEN s_14_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_13(183) WHEN s_14_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_13(184) WHEN s_14_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_13(185) WHEN s_14_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_13(186) WHEN s_14_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_13(187) WHEN s_14_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_13(188) WHEN s_14_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_13(189) WHEN s_14_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_13(190) WHEN s_14_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_13(191) WHEN s_14_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_13(192) WHEN s_14_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_13(193) WHEN s_14_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_13(194) WHEN s_14_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_13(195) WHEN s_14_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_13(196) WHEN s_14_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_13(197) WHEN s_14_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_13(198) WHEN s_14_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_13(199) WHEN s_14_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_13(200) WHEN s_14_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_13(201) WHEN s_14_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_13(202) WHEN s_14_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_13(203) WHEN s_14_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_13(204) WHEN s_14_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_13(205) WHEN s_14_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_13(206) WHEN s_14_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_13(207) WHEN s_14_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_13(208) WHEN s_14_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_13(209) WHEN s_14_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_13(210) WHEN s_14_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_13(211) WHEN s_14_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_13(212) WHEN s_14_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_13(213) WHEN s_14_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_13(214) WHEN s_14_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_13(215) WHEN s_14_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_13(216) WHEN s_14_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_13(217) WHEN s_14_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_13(218) WHEN s_14_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_13(219) WHEN s_14_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_13(220) WHEN s_14_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_13(221) WHEN s_14_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_13(222) WHEN s_14_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_13(223) WHEN s_14_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_13(224) WHEN s_14_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_13(225) WHEN s_14_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_13(226) WHEN s_14_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_13(227) WHEN s_14_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_13(228) WHEN s_14_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_13(229) WHEN s_14_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_13(230) WHEN s_14_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_13(231) WHEN s_14_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_13(232) WHEN s_14_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_13(233) WHEN s_14_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_13(234) WHEN s_14_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_13(235) WHEN s_14_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_13(236) WHEN s_14_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_13(237) WHEN s_14_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_13(238) WHEN s_14_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_13(239) WHEN s_14_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_13(240) WHEN s_14_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_13(241) WHEN s_14_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_13(242) WHEN s_14_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_13(243) WHEN s_14_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_13(244) WHEN s_14_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_13(245) WHEN s_14_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_13(246) WHEN s_14_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_13(247) WHEN s_14_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_13(248) WHEN s_14_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_13(249) WHEN s_14_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_13(250) WHEN s_14_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_13(251) WHEN s_14_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_13(252) WHEN s_14_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_13(253) WHEN s_14_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_13(254) WHEN s_14_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_13(255);

  
  out0_136 <= gmul2_13(0) WHEN s_13_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_13(1) WHEN s_13_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_13(2) WHEN s_13_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_13(3) WHEN s_13_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_13(4) WHEN s_13_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_13(5) WHEN s_13_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_13(6) WHEN s_13_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_13(7) WHEN s_13_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_13(8) WHEN s_13_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_13(9) WHEN s_13_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_13(10) WHEN s_13_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_13(11) WHEN s_13_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_13(12) WHEN s_13_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_13(13) WHEN s_13_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_13(14) WHEN s_13_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_13(15) WHEN s_13_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_13(16) WHEN s_13_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_13(17) WHEN s_13_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_13(18) WHEN s_13_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_13(19) WHEN s_13_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_13(20) WHEN s_13_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_13(21) WHEN s_13_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_13(22) WHEN s_13_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_13(23) WHEN s_13_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_13(24) WHEN s_13_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_13(25) WHEN s_13_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_13(26) WHEN s_13_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_13(27) WHEN s_13_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_13(28) WHEN s_13_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_13(29) WHEN s_13_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_13(30) WHEN s_13_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_13(31) WHEN s_13_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_13(32) WHEN s_13_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_13(33) WHEN s_13_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_13(34) WHEN s_13_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_13(35) WHEN s_13_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_13(36) WHEN s_13_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_13(37) WHEN s_13_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_13(38) WHEN s_13_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_13(39) WHEN s_13_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_13(40) WHEN s_13_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_13(41) WHEN s_13_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_13(42) WHEN s_13_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_13(43) WHEN s_13_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_13(44) WHEN s_13_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_13(45) WHEN s_13_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_13(46) WHEN s_13_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_13(47) WHEN s_13_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_13(48) WHEN s_13_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_13(49) WHEN s_13_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_13(50) WHEN s_13_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_13(51) WHEN s_13_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_13(52) WHEN s_13_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_13(53) WHEN s_13_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_13(54) WHEN s_13_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_13(55) WHEN s_13_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_13(56) WHEN s_13_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_13(57) WHEN s_13_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_13(58) WHEN s_13_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_13(59) WHEN s_13_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_13(60) WHEN s_13_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_13(61) WHEN s_13_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_13(62) WHEN s_13_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_13(63) WHEN s_13_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_13(64) WHEN s_13_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_13(65) WHEN s_13_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_13(66) WHEN s_13_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_13(67) WHEN s_13_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_13(68) WHEN s_13_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_13(69) WHEN s_13_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_13(70) WHEN s_13_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_13(71) WHEN s_13_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_13(72) WHEN s_13_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_13(73) WHEN s_13_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_13(74) WHEN s_13_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_13(75) WHEN s_13_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_13(76) WHEN s_13_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_13(77) WHEN s_13_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_13(78) WHEN s_13_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_13(79) WHEN s_13_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_13(80) WHEN s_13_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_13(81) WHEN s_13_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_13(82) WHEN s_13_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_13(83) WHEN s_13_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_13(84) WHEN s_13_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_13(85) WHEN s_13_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_13(86) WHEN s_13_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_13(87) WHEN s_13_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_13(88) WHEN s_13_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_13(89) WHEN s_13_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_13(90) WHEN s_13_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_13(91) WHEN s_13_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_13(92) WHEN s_13_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_13(93) WHEN s_13_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_13(94) WHEN s_13_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_13(95) WHEN s_13_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_13(96) WHEN s_13_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_13(97) WHEN s_13_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_13(98) WHEN s_13_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_13(99) WHEN s_13_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_13(100) WHEN s_13_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_13(101) WHEN s_13_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_13(102) WHEN s_13_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_13(103) WHEN s_13_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_13(104) WHEN s_13_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_13(105) WHEN s_13_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_13(106) WHEN s_13_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_13(107) WHEN s_13_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_13(108) WHEN s_13_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_13(109) WHEN s_13_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_13(110) WHEN s_13_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_13(111) WHEN s_13_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_13(112) WHEN s_13_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_13(113) WHEN s_13_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_13(114) WHEN s_13_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_13(115) WHEN s_13_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_13(116) WHEN s_13_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_13(117) WHEN s_13_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_13(118) WHEN s_13_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_13(119) WHEN s_13_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_13(120) WHEN s_13_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_13(121) WHEN s_13_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_13(122) WHEN s_13_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_13(123) WHEN s_13_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_13(124) WHEN s_13_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_13(125) WHEN s_13_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_13(126) WHEN s_13_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_13(127) WHEN s_13_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_13(128) WHEN s_13_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_13(129) WHEN s_13_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_13(130) WHEN s_13_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_13(131) WHEN s_13_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_13(132) WHEN s_13_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_13(133) WHEN s_13_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_13(134) WHEN s_13_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_13(135) WHEN s_13_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_13(136) WHEN s_13_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_13(137) WHEN s_13_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_13(138) WHEN s_13_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_13(139) WHEN s_13_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_13(140) WHEN s_13_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_13(141) WHEN s_13_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_13(142) WHEN s_13_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_13(143) WHEN s_13_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_13(144) WHEN s_13_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_13(145) WHEN s_13_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_13(146) WHEN s_13_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_13(147) WHEN s_13_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_13(148) WHEN s_13_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_13(149) WHEN s_13_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_13(150) WHEN s_13_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_13(151) WHEN s_13_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_13(152) WHEN s_13_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_13(153) WHEN s_13_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_13(154) WHEN s_13_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_13(155) WHEN s_13_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_13(156) WHEN s_13_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_13(157) WHEN s_13_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_13(158) WHEN s_13_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_13(159) WHEN s_13_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_13(160) WHEN s_13_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_13(161) WHEN s_13_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_13(162) WHEN s_13_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_13(163) WHEN s_13_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_13(164) WHEN s_13_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_13(165) WHEN s_13_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_13(166) WHEN s_13_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_13(167) WHEN s_13_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_13(168) WHEN s_13_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_13(169) WHEN s_13_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_13(170) WHEN s_13_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_13(171) WHEN s_13_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_13(172) WHEN s_13_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_13(173) WHEN s_13_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_13(174) WHEN s_13_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_13(175) WHEN s_13_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_13(176) WHEN s_13_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_13(177) WHEN s_13_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_13(178) WHEN s_13_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_13(179) WHEN s_13_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_13(180) WHEN s_13_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_13(181) WHEN s_13_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_13(182) WHEN s_13_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_13(183) WHEN s_13_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_13(184) WHEN s_13_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_13(185) WHEN s_13_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_13(186) WHEN s_13_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_13(187) WHEN s_13_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_13(188) WHEN s_13_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_13(189) WHEN s_13_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_13(190) WHEN s_13_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_13(191) WHEN s_13_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_13(192) WHEN s_13_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_13(193) WHEN s_13_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_13(194) WHEN s_13_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_13(195) WHEN s_13_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_13(196) WHEN s_13_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_13(197) WHEN s_13_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_13(198) WHEN s_13_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_13(199) WHEN s_13_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_13(200) WHEN s_13_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_13(201) WHEN s_13_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_13(202) WHEN s_13_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_13(203) WHEN s_13_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_13(204) WHEN s_13_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_13(205) WHEN s_13_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_13(206) WHEN s_13_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_13(207) WHEN s_13_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_13(208) WHEN s_13_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_13(209) WHEN s_13_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_13(210) WHEN s_13_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_13(211) WHEN s_13_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_13(212) WHEN s_13_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_13(213) WHEN s_13_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_13(214) WHEN s_13_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_13(215) WHEN s_13_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_13(216) WHEN s_13_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_13(217) WHEN s_13_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_13(218) WHEN s_13_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_13(219) WHEN s_13_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_13(220) WHEN s_13_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_13(221) WHEN s_13_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_13(222) WHEN s_13_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_13(223) WHEN s_13_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_13(224) WHEN s_13_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_13(225) WHEN s_13_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_13(226) WHEN s_13_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_13(227) WHEN s_13_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_13(228) WHEN s_13_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_13(229) WHEN s_13_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_13(230) WHEN s_13_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_13(231) WHEN s_13_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_13(232) WHEN s_13_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_13(233) WHEN s_13_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_13(234) WHEN s_13_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_13(235) WHEN s_13_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_13(236) WHEN s_13_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_13(237) WHEN s_13_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_13(238) WHEN s_13_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_13(239) WHEN s_13_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_13(240) WHEN s_13_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_13(241) WHEN s_13_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_13(242) WHEN s_13_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_13(243) WHEN s_13_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_13(244) WHEN s_13_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_13(245) WHEN s_13_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_13(246) WHEN s_13_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_13(247) WHEN s_13_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_13(248) WHEN s_13_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_13(249) WHEN s_13_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_13(250) WHEN s_13_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_13(251) WHEN s_13_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_13(252) WHEN s_13_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_13(253) WHEN s_13_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_13(254) WHEN s_13_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_13(255);

  out0_137 <= s_12_1 XOR out0_136;

  b2 <= out0_137 XOR out0_135;

  out0_138 <= b2 XOR s_15_1;

  s_15_1 <= s_s_4(15);

  s_14_1 <= s_s_4(14);

  s_13_1 <= s_s_4(13);

  
  out0_139 <= gmul3_12(0) WHEN s_13_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_12(1) WHEN s_13_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_12(2) WHEN s_13_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_12(3) WHEN s_13_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_12(4) WHEN s_13_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_12(5) WHEN s_13_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_12(6) WHEN s_13_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_12(7) WHEN s_13_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_12(8) WHEN s_13_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_12(9) WHEN s_13_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_12(10) WHEN s_13_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_12(11) WHEN s_13_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_12(12) WHEN s_13_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_12(13) WHEN s_13_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_12(14) WHEN s_13_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_12(15) WHEN s_13_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_12(16) WHEN s_13_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_12(17) WHEN s_13_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_12(18) WHEN s_13_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_12(19) WHEN s_13_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_12(20) WHEN s_13_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_12(21) WHEN s_13_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_12(22) WHEN s_13_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_12(23) WHEN s_13_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_12(24) WHEN s_13_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_12(25) WHEN s_13_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_12(26) WHEN s_13_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_12(27) WHEN s_13_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_12(28) WHEN s_13_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_12(29) WHEN s_13_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_12(30) WHEN s_13_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_12(31) WHEN s_13_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_12(32) WHEN s_13_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_12(33) WHEN s_13_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_12(34) WHEN s_13_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_12(35) WHEN s_13_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_12(36) WHEN s_13_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_12(37) WHEN s_13_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_12(38) WHEN s_13_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_12(39) WHEN s_13_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_12(40) WHEN s_13_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_12(41) WHEN s_13_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_12(42) WHEN s_13_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_12(43) WHEN s_13_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_12(44) WHEN s_13_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_12(45) WHEN s_13_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_12(46) WHEN s_13_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_12(47) WHEN s_13_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_12(48) WHEN s_13_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_12(49) WHEN s_13_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_12(50) WHEN s_13_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_12(51) WHEN s_13_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_12(52) WHEN s_13_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_12(53) WHEN s_13_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_12(54) WHEN s_13_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_12(55) WHEN s_13_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_12(56) WHEN s_13_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_12(57) WHEN s_13_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_12(58) WHEN s_13_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_12(59) WHEN s_13_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_12(60) WHEN s_13_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_12(61) WHEN s_13_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_12(62) WHEN s_13_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_12(63) WHEN s_13_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_12(64) WHEN s_13_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_12(65) WHEN s_13_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_12(66) WHEN s_13_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_12(67) WHEN s_13_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_12(68) WHEN s_13_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_12(69) WHEN s_13_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_12(70) WHEN s_13_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_12(71) WHEN s_13_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_12(72) WHEN s_13_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_12(73) WHEN s_13_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_12(74) WHEN s_13_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_12(75) WHEN s_13_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_12(76) WHEN s_13_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_12(77) WHEN s_13_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_12(78) WHEN s_13_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_12(79) WHEN s_13_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_12(80) WHEN s_13_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_12(81) WHEN s_13_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_12(82) WHEN s_13_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_12(83) WHEN s_13_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_12(84) WHEN s_13_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_12(85) WHEN s_13_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_12(86) WHEN s_13_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_12(87) WHEN s_13_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_12(88) WHEN s_13_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_12(89) WHEN s_13_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_12(90) WHEN s_13_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_12(91) WHEN s_13_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_12(92) WHEN s_13_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_12(93) WHEN s_13_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_12(94) WHEN s_13_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_12(95) WHEN s_13_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_12(96) WHEN s_13_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_12(97) WHEN s_13_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_12(98) WHEN s_13_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_12(99) WHEN s_13_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_12(100) WHEN s_13_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_12(101) WHEN s_13_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_12(102) WHEN s_13_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_12(103) WHEN s_13_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_12(104) WHEN s_13_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_12(105) WHEN s_13_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_12(106) WHEN s_13_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_12(107) WHEN s_13_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_12(108) WHEN s_13_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_12(109) WHEN s_13_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_12(110) WHEN s_13_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_12(111) WHEN s_13_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_12(112) WHEN s_13_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_12(113) WHEN s_13_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_12(114) WHEN s_13_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_12(115) WHEN s_13_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_12(116) WHEN s_13_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_12(117) WHEN s_13_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_12(118) WHEN s_13_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_12(119) WHEN s_13_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_12(120) WHEN s_13_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_12(121) WHEN s_13_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_12(122) WHEN s_13_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_12(123) WHEN s_13_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_12(124) WHEN s_13_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_12(125) WHEN s_13_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_12(126) WHEN s_13_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_12(127) WHEN s_13_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_12(128) WHEN s_13_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_12(129) WHEN s_13_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_12(130) WHEN s_13_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_12(131) WHEN s_13_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_12(132) WHEN s_13_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_12(133) WHEN s_13_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_12(134) WHEN s_13_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_12(135) WHEN s_13_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_12(136) WHEN s_13_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_12(137) WHEN s_13_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_12(138) WHEN s_13_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_12(139) WHEN s_13_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_12(140) WHEN s_13_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_12(141) WHEN s_13_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_12(142) WHEN s_13_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_12(143) WHEN s_13_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_12(144) WHEN s_13_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_12(145) WHEN s_13_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_12(146) WHEN s_13_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_12(147) WHEN s_13_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_12(148) WHEN s_13_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_12(149) WHEN s_13_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_12(150) WHEN s_13_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_12(151) WHEN s_13_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_12(152) WHEN s_13_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_12(153) WHEN s_13_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_12(154) WHEN s_13_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_12(155) WHEN s_13_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_12(156) WHEN s_13_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_12(157) WHEN s_13_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_12(158) WHEN s_13_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_12(159) WHEN s_13_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_12(160) WHEN s_13_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_12(161) WHEN s_13_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_12(162) WHEN s_13_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_12(163) WHEN s_13_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_12(164) WHEN s_13_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_12(165) WHEN s_13_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_12(166) WHEN s_13_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_12(167) WHEN s_13_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_12(168) WHEN s_13_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_12(169) WHEN s_13_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_12(170) WHEN s_13_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_12(171) WHEN s_13_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_12(172) WHEN s_13_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_12(173) WHEN s_13_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_12(174) WHEN s_13_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_12(175) WHEN s_13_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_12(176) WHEN s_13_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_12(177) WHEN s_13_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_12(178) WHEN s_13_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_12(179) WHEN s_13_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_12(180) WHEN s_13_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_12(181) WHEN s_13_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_12(182) WHEN s_13_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_12(183) WHEN s_13_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_12(184) WHEN s_13_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_12(185) WHEN s_13_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_12(186) WHEN s_13_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_12(187) WHEN s_13_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_12(188) WHEN s_13_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_12(189) WHEN s_13_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_12(190) WHEN s_13_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_12(191) WHEN s_13_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_12(192) WHEN s_13_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_12(193) WHEN s_13_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_12(194) WHEN s_13_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_12(195) WHEN s_13_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_12(196) WHEN s_13_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_12(197) WHEN s_13_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_12(198) WHEN s_13_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_12(199) WHEN s_13_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_12(200) WHEN s_13_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_12(201) WHEN s_13_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_12(202) WHEN s_13_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_12(203) WHEN s_13_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_12(204) WHEN s_13_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_12(205) WHEN s_13_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_12(206) WHEN s_13_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_12(207) WHEN s_13_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_12(208) WHEN s_13_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_12(209) WHEN s_13_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_12(210) WHEN s_13_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_12(211) WHEN s_13_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_12(212) WHEN s_13_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_12(213) WHEN s_13_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_12(214) WHEN s_13_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_12(215) WHEN s_13_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_12(216) WHEN s_13_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_12(217) WHEN s_13_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_12(218) WHEN s_13_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_12(219) WHEN s_13_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_12(220) WHEN s_13_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_12(221) WHEN s_13_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_12(222) WHEN s_13_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_12(223) WHEN s_13_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_12(224) WHEN s_13_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_12(225) WHEN s_13_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_12(226) WHEN s_13_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_12(227) WHEN s_13_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_12(228) WHEN s_13_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_12(229) WHEN s_13_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_12(230) WHEN s_13_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_12(231) WHEN s_13_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_12(232) WHEN s_13_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_12(233) WHEN s_13_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_12(234) WHEN s_13_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_12(235) WHEN s_13_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_12(236) WHEN s_13_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_12(237) WHEN s_13_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_12(238) WHEN s_13_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_12(239) WHEN s_13_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_12(240) WHEN s_13_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_12(241) WHEN s_13_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_12(242) WHEN s_13_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_12(243) WHEN s_13_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_12(244) WHEN s_13_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_12(245) WHEN s_13_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_12(246) WHEN s_13_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_12(247) WHEN s_13_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_12(248) WHEN s_13_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_12(249) WHEN s_13_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_12(250) WHEN s_13_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_12(251) WHEN s_13_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_12(252) WHEN s_13_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_12(253) WHEN s_13_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_12(254) WHEN s_13_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_12(255);

  s_12_1 <= s_s_4(12);

  
  out0_140 <= gmul2_12(0) WHEN s_12_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_12(1) WHEN s_12_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_12(2) WHEN s_12_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_12(3) WHEN s_12_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_12(4) WHEN s_12_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_12(5) WHEN s_12_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_12(6) WHEN s_12_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_12(7) WHEN s_12_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_12(8) WHEN s_12_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_12(9) WHEN s_12_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_12(10) WHEN s_12_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_12(11) WHEN s_12_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_12(12) WHEN s_12_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_12(13) WHEN s_12_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_12(14) WHEN s_12_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_12(15) WHEN s_12_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_12(16) WHEN s_12_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_12(17) WHEN s_12_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_12(18) WHEN s_12_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_12(19) WHEN s_12_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_12(20) WHEN s_12_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_12(21) WHEN s_12_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_12(22) WHEN s_12_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_12(23) WHEN s_12_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_12(24) WHEN s_12_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_12(25) WHEN s_12_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_12(26) WHEN s_12_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_12(27) WHEN s_12_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_12(28) WHEN s_12_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_12(29) WHEN s_12_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_12(30) WHEN s_12_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_12(31) WHEN s_12_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_12(32) WHEN s_12_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_12(33) WHEN s_12_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_12(34) WHEN s_12_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_12(35) WHEN s_12_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_12(36) WHEN s_12_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_12(37) WHEN s_12_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_12(38) WHEN s_12_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_12(39) WHEN s_12_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_12(40) WHEN s_12_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_12(41) WHEN s_12_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_12(42) WHEN s_12_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_12(43) WHEN s_12_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_12(44) WHEN s_12_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_12(45) WHEN s_12_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_12(46) WHEN s_12_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_12(47) WHEN s_12_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_12(48) WHEN s_12_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_12(49) WHEN s_12_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_12(50) WHEN s_12_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_12(51) WHEN s_12_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_12(52) WHEN s_12_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_12(53) WHEN s_12_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_12(54) WHEN s_12_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_12(55) WHEN s_12_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_12(56) WHEN s_12_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_12(57) WHEN s_12_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_12(58) WHEN s_12_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_12(59) WHEN s_12_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_12(60) WHEN s_12_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_12(61) WHEN s_12_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_12(62) WHEN s_12_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_12(63) WHEN s_12_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_12(64) WHEN s_12_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_12(65) WHEN s_12_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_12(66) WHEN s_12_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_12(67) WHEN s_12_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_12(68) WHEN s_12_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_12(69) WHEN s_12_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_12(70) WHEN s_12_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_12(71) WHEN s_12_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_12(72) WHEN s_12_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_12(73) WHEN s_12_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_12(74) WHEN s_12_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_12(75) WHEN s_12_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_12(76) WHEN s_12_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_12(77) WHEN s_12_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_12(78) WHEN s_12_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_12(79) WHEN s_12_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_12(80) WHEN s_12_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_12(81) WHEN s_12_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_12(82) WHEN s_12_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_12(83) WHEN s_12_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_12(84) WHEN s_12_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_12(85) WHEN s_12_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_12(86) WHEN s_12_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_12(87) WHEN s_12_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_12(88) WHEN s_12_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_12(89) WHEN s_12_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_12(90) WHEN s_12_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_12(91) WHEN s_12_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_12(92) WHEN s_12_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_12(93) WHEN s_12_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_12(94) WHEN s_12_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_12(95) WHEN s_12_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_12(96) WHEN s_12_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_12(97) WHEN s_12_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_12(98) WHEN s_12_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_12(99) WHEN s_12_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_12(100) WHEN s_12_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_12(101) WHEN s_12_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_12(102) WHEN s_12_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_12(103) WHEN s_12_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_12(104) WHEN s_12_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_12(105) WHEN s_12_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_12(106) WHEN s_12_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_12(107) WHEN s_12_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_12(108) WHEN s_12_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_12(109) WHEN s_12_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_12(110) WHEN s_12_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_12(111) WHEN s_12_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_12(112) WHEN s_12_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_12(113) WHEN s_12_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_12(114) WHEN s_12_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_12(115) WHEN s_12_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_12(116) WHEN s_12_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_12(117) WHEN s_12_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_12(118) WHEN s_12_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_12(119) WHEN s_12_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_12(120) WHEN s_12_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_12(121) WHEN s_12_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_12(122) WHEN s_12_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_12(123) WHEN s_12_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_12(124) WHEN s_12_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_12(125) WHEN s_12_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_12(126) WHEN s_12_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_12(127) WHEN s_12_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_12(128) WHEN s_12_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_12(129) WHEN s_12_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_12(130) WHEN s_12_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_12(131) WHEN s_12_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_12(132) WHEN s_12_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_12(133) WHEN s_12_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_12(134) WHEN s_12_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_12(135) WHEN s_12_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_12(136) WHEN s_12_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_12(137) WHEN s_12_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_12(138) WHEN s_12_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_12(139) WHEN s_12_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_12(140) WHEN s_12_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_12(141) WHEN s_12_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_12(142) WHEN s_12_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_12(143) WHEN s_12_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_12(144) WHEN s_12_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_12(145) WHEN s_12_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_12(146) WHEN s_12_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_12(147) WHEN s_12_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_12(148) WHEN s_12_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_12(149) WHEN s_12_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_12(150) WHEN s_12_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_12(151) WHEN s_12_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_12(152) WHEN s_12_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_12(153) WHEN s_12_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_12(154) WHEN s_12_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_12(155) WHEN s_12_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_12(156) WHEN s_12_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_12(157) WHEN s_12_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_12(158) WHEN s_12_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_12(159) WHEN s_12_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_12(160) WHEN s_12_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_12(161) WHEN s_12_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_12(162) WHEN s_12_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_12(163) WHEN s_12_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_12(164) WHEN s_12_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_12(165) WHEN s_12_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_12(166) WHEN s_12_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_12(167) WHEN s_12_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_12(168) WHEN s_12_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_12(169) WHEN s_12_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_12(170) WHEN s_12_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_12(171) WHEN s_12_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_12(172) WHEN s_12_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_12(173) WHEN s_12_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_12(174) WHEN s_12_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_12(175) WHEN s_12_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_12(176) WHEN s_12_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_12(177) WHEN s_12_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_12(178) WHEN s_12_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_12(179) WHEN s_12_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_12(180) WHEN s_12_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_12(181) WHEN s_12_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_12(182) WHEN s_12_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_12(183) WHEN s_12_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_12(184) WHEN s_12_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_12(185) WHEN s_12_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_12(186) WHEN s_12_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_12(187) WHEN s_12_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_12(188) WHEN s_12_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_12(189) WHEN s_12_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_12(190) WHEN s_12_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_12(191) WHEN s_12_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_12(192) WHEN s_12_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_12(193) WHEN s_12_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_12(194) WHEN s_12_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_12(195) WHEN s_12_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_12(196) WHEN s_12_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_12(197) WHEN s_12_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_12(198) WHEN s_12_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_12(199) WHEN s_12_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_12(200) WHEN s_12_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_12(201) WHEN s_12_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_12(202) WHEN s_12_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_12(203) WHEN s_12_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_12(204) WHEN s_12_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_12(205) WHEN s_12_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_12(206) WHEN s_12_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_12(207) WHEN s_12_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_12(208) WHEN s_12_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_12(209) WHEN s_12_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_12(210) WHEN s_12_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_12(211) WHEN s_12_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_12(212) WHEN s_12_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_12(213) WHEN s_12_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_12(214) WHEN s_12_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_12(215) WHEN s_12_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_12(216) WHEN s_12_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_12(217) WHEN s_12_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_12(218) WHEN s_12_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_12(219) WHEN s_12_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_12(220) WHEN s_12_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_12(221) WHEN s_12_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_12(222) WHEN s_12_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_12(223) WHEN s_12_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_12(224) WHEN s_12_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_12(225) WHEN s_12_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_12(226) WHEN s_12_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_12(227) WHEN s_12_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_12(228) WHEN s_12_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_12(229) WHEN s_12_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_12(230) WHEN s_12_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_12(231) WHEN s_12_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_12(232) WHEN s_12_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_12(233) WHEN s_12_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_12(234) WHEN s_12_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_12(235) WHEN s_12_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_12(236) WHEN s_12_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_12(237) WHEN s_12_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_12(238) WHEN s_12_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_12(239) WHEN s_12_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_12(240) WHEN s_12_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_12(241) WHEN s_12_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_12(242) WHEN s_12_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_12(243) WHEN s_12_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_12(244) WHEN s_12_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_12(245) WHEN s_12_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_12(246) WHEN s_12_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_12(247) WHEN s_12_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_12(248) WHEN s_12_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_12(249) WHEN s_12_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_12(250) WHEN s_12_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_12(251) WHEN s_12_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_12(252) WHEN s_12_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_12(253) WHEN s_12_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_12(254) WHEN s_12_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_12(255);

  out0_141 <= out0_140 XOR out0_139;

  b1 <= out0_141 XOR s_14_1;

  out0_142 <= b1 XOR s_15_1;

  
  out0_143 <= gmul2_11(0) WHEN s_11_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_11(1) WHEN s_11_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_11(2) WHEN s_11_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_11(3) WHEN s_11_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_11(4) WHEN s_11_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_11(5) WHEN s_11_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_11(6) WHEN s_11_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_11(7) WHEN s_11_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_11(8) WHEN s_11_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_11(9) WHEN s_11_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_11(10) WHEN s_11_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_11(11) WHEN s_11_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_11(12) WHEN s_11_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_11(13) WHEN s_11_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_11(14) WHEN s_11_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_11(15) WHEN s_11_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_11(16) WHEN s_11_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_11(17) WHEN s_11_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_11(18) WHEN s_11_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_11(19) WHEN s_11_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_11(20) WHEN s_11_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_11(21) WHEN s_11_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_11(22) WHEN s_11_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_11(23) WHEN s_11_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_11(24) WHEN s_11_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_11(25) WHEN s_11_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_11(26) WHEN s_11_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_11(27) WHEN s_11_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_11(28) WHEN s_11_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_11(29) WHEN s_11_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_11(30) WHEN s_11_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_11(31) WHEN s_11_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_11(32) WHEN s_11_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_11(33) WHEN s_11_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_11(34) WHEN s_11_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_11(35) WHEN s_11_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_11(36) WHEN s_11_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_11(37) WHEN s_11_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_11(38) WHEN s_11_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_11(39) WHEN s_11_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_11(40) WHEN s_11_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_11(41) WHEN s_11_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_11(42) WHEN s_11_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_11(43) WHEN s_11_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_11(44) WHEN s_11_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_11(45) WHEN s_11_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_11(46) WHEN s_11_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_11(47) WHEN s_11_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_11(48) WHEN s_11_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_11(49) WHEN s_11_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_11(50) WHEN s_11_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_11(51) WHEN s_11_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_11(52) WHEN s_11_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_11(53) WHEN s_11_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_11(54) WHEN s_11_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_11(55) WHEN s_11_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_11(56) WHEN s_11_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_11(57) WHEN s_11_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_11(58) WHEN s_11_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_11(59) WHEN s_11_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_11(60) WHEN s_11_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_11(61) WHEN s_11_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_11(62) WHEN s_11_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_11(63) WHEN s_11_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_11(64) WHEN s_11_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_11(65) WHEN s_11_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_11(66) WHEN s_11_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_11(67) WHEN s_11_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_11(68) WHEN s_11_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_11(69) WHEN s_11_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_11(70) WHEN s_11_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_11(71) WHEN s_11_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_11(72) WHEN s_11_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_11(73) WHEN s_11_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_11(74) WHEN s_11_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_11(75) WHEN s_11_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_11(76) WHEN s_11_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_11(77) WHEN s_11_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_11(78) WHEN s_11_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_11(79) WHEN s_11_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_11(80) WHEN s_11_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_11(81) WHEN s_11_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_11(82) WHEN s_11_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_11(83) WHEN s_11_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_11(84) WHEN s_11_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_11(85) WHEN s_11_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_11(86) WHEN s_11_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_11(87) WHEN s_11_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_11(88) WHEN s_11_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_11(89) WHEN s_11_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_11(90) WHEN s_11_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_11(91) WHEN s_11_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_11(92) WHEN s_11_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_11(93) WHEN s_11_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_11(94) WHEN s_11_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_11(95) WHEN s_11_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_11(96) WHEN s_11_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_11(97) WHEN s_11_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_11(98) WHEN s_11_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_11(99) WHEN s_11_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_11(100) WHEN s_11_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_11(101) WHEN s_11_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_11(102) WHEN s_11_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_11(103) WHEN s_11_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_11(104) WHEN s_11_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_11(105) WHEN s_11_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_11(106) WHEN s_11_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_11(107) WHEN s_11_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_11(108) WHEN s_11_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_11(109) WHEN s_11_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_11(110) WHEN s_11_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_11(111) WHEN s_11_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_11(112) WHEN s_11_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_11(113) WHEN s_11_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_11(114) WHEN s_11_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_11(115) WHEN s_11_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_11(116) WHEN s_11_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_11(117) WHEN s_11_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_11(118) WHEN s_11_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_11(119) WHEN s_11_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_11(120) WHEN s_11_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_11(121) WHEN s_11_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_11(122) WHEN s_11_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_11(123) WHEN s_11_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_11(124) WHEN s_11_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_11(125) WHEN s_11_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_11(126) WHEN s_11_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_11(127) WHEN s_11_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_11(128) WHEN s_11_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_11(129) WHEN s_11_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_11(130) WHEN s_11_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_11(131) WHEN s_11_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_11(132) WHEN s_11_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_11(133) WHEN s_11_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_11(134) WHEN s_11_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_11(135) WHEN s_11_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_11(136) WHEN s_11_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_11(137) WHEN s_11_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_11(138) WHEN s_11_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_11(139) WHEN s_11_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_11(140) WHEN s_11_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_11(141) WHEN s_11_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_11(142) WHEN s_11_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_11(143) WHEN s_11_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_11(144) WHEN s_11_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_11(145) WHEN s_11_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_11(146) WHEN s_11_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_11(147) WHEN s_11_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_11(148) WHEN s_11_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_11(149) WHEN s_11_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_11(150) WHEN s_11_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_11(151) WHEN s_11_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_11(152) WHEN s_11_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_11(153) WHEN s_11_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_11(154) WHEN s_11_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_11(155) WHEN s_11_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_11(156) WHEN s_11_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_11(157) WHEN s_11_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_11(158) WHEN s_11_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_11(159) WHEN s_11_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_11(160) WHEN s_11_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_11(161) WHEN s_11_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_11(162) WHEN s_11_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_11(163) WHEN s_11_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_11(164) WHEN s_11_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_11(165) WHEN s_11_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_11(166) WHEN s_11_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_11(167) WHEN s_11_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_11(168) WHEN s_11_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_11(169) WHEN s_11_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_11(170) WHEN s_11_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_11(171) WHEN s_11_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_11(172) WHEN s_11_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_11(173) WHEN s_11_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_11(174) WHEN s_11_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_11(175) WHEN s_11_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_11(176) WHEN s_11_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_11(177) WHEN s_11_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_11(178) WHEN s_11_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_11(179) WHEN s_11_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_11(180) WHEN s_11_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_11(181) WHEN s_11_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_11(182) WHEN s_11_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_11(183) WHEN s_11_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_11(184) WHEN s_11_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_11(185) WHEN s_11_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_11(186) WHEN s_11_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_11(187) WHEN s_11_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_11(188) WHEN s_11_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_11(189) WHEN s_11_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_11(190) WHEN s_11_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_11(191) WHEN s_11_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_11(192) WHEN s_11_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_11(193) WHEN s_11_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_11(194) WHEN s_11_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_11(195) WHEN s_11_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_11(196) WHEN s_11_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_11(197) WHEN s_11_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_11(198) WHEN s_11_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_11(199) WHEN s_11_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_11(200) WHEN s_11_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_11(201) WHEN s_11_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_11(202) WHEN s_11_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_11(203) WHEN s_11_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_11(204) WHEN s_11_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_11(205) WHEN s_11_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_11(206) WHEN s_11_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_11(207) WHEN s_11_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_11(208) WHEN s_11_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_11(209) WHEN s_11_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_11(210) WHEN s_11_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_11(211) WHEN s_11_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_11(212) WHEN s_11_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_11(213) WHEN s_11_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_11(214) WHEN s_11_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_11(215) WHEN s_11_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_11(216) WHEN s_11_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_11(217) WHEN s_11_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_11(218) WHEN s_11_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_11(219) WHEN s_11_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_11(220) WHEN s_11_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_11(221) WHEN s_11_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_11(222) WHEN s_11_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_11(223) WHEN s_11_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_11(224) WHEN s_11_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_11(225) WHEN s_11_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_11(226) WHEN s_11_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_11(227) WHEN s_11_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_11(228) WHEN s_11_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_11(229) WHEN s_11_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_11(230) WHEN s_11_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_11(231) WHEN s_11_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_11(232) WHEN s_11_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_11(233) WHEN s_11_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_11(234) WHEN s_11_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_11(235) WHEN s_11_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_11(236) WHEN s_11_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_11(237) WHEN s_11_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_11(238) WHEN s_11_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_11(239) WHEN s_11_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_11(240) WHEN s_11_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_11(241) WHEN s_11_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_11(242) WHEN s_11_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_11(243) WHEN s_11_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_11(244) WHEN s_11_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_11(245) WHEN s_11_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_11(246) WHEN s_11_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_11(247) WHEN s_11_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_11(248) WHEN s_11_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_11(249) WHEN s_11_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_11(250) WHEN s_11_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_11(251) WHEN s_11_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_11(252) WHEN s_11_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_11(253) WHEN s_11_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_11(254) WHEN s_11_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_11(255);

  
  out0_144 <= gmul3_11(0) WHEN s_8_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_11(1) WHEN s_8_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_11(2) WHEN s_8_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_11(3) WHEN s_8_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_11(4) WHEN s_8_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_11(5) WHEN s_8_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_11(6) WHEN s_8_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_11(7) WHEN s_8_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_11(8) WHEN s_8_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_11(9) WHEN s_8_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_11(10) WHEN s_8_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_11(11) WHEN s_8_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_11(12) WHEN s_8_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_11(13) WHEN s_8_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_11(14) WHEN s_8_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_11(15) WHEN s_8_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_11(16) WHEN s_8_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_11(17) WHEN s_8_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_11(18) WHEN s_8_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_11(19) WHEN s_8_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_11(20) WHEN s_8_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_11(21) WHEN s_8_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_11(22) WHEN s_8_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_11(23) WHEN s_8_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_11(24) WHEN s_8_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_11(25) WHEN s_8_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_11(26) WHEN s_8_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_11(27) WHEN s_8_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_11(28) WHEN s_8_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_11(29) WHEN s_8_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_11(30) WHEN s_8_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_11(31) WHEN s_8_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_11(32) WHEN s_8_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_11(33) WHEN s_8_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_11(34) WHEN s_8_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_11(35) WHEN s_8_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_11(36) WHEN s_8_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_11(37) WHEN s_8_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_11(38) WHEN s_8_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_11(39) WHEN s_8_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_11(40) WHEN s_8_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_11(41) WHEN s_8_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_11(42) WHEN s_8_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_11(43) WHEN s_8_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_11(44) WHEN s_8_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_11(45) WHEN s_8_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_11(46) WHEN s_8_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_11(47) WHEN s_8_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_11(48) WHEN s_8_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_11(49) WHEN s_8_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_11(50) WHEN s_8_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_11(51) WHEN s_8_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_11(52) WHEN s_8_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_11(53) WHEN s_8_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_11(54) WHEN s_8_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_11(55) WHEN s_8_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_11(56) WHEN s_8_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_11(57) WHEN s_8_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_11(58) WHEN s_8_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_11(59) WHEN s_8_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_11(60) WHEN s_8_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_11(61) WHEN s_8_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_11(62) WHEN s_8_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_11(63) WHEN s_8_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_11(64) WHEN s_8_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_11(65) WHEN s_8_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_11(66) WHEN s_8_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_11(67) WHEN s_8_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_11(68) WHEN s_8_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_11(69) WHEN s_8_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_11(70) WHEN s_8_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_11(71) WHEN s_8_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_11(72) WHEN s_8_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_11(73) WHEN s_8_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_11(74) WHEN s_8_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_11(75) WHEN s_8_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_11(76) WHEN s_8_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_11(77) WHEN s_8_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_11(78) WHEN s_8_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_11(79) WHEN s_8_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_11(80) WHEN s_8_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_11(81) WHEN s_8_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_11(82) WHEN s_8_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_11(83) WHEN s_8_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_11(84) WHEN s_8_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_11(85) WHEN s_8_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_11(86) WHEN s_8_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_11(87) WHEN s_8_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_11(88) WHEN s_8_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_11(89) WHEN s_8_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_11(90) WHEN s_8_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_11(91) WHEN s_8_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_11(92) WHEN s_8_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_11(93) WHEN s_8_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_11(94) WHEN s_8_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_11(95) WHEN s_8_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_11(96) WHEN s_8_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_11(97) WHEN s_8_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_11(98) WHEN s_8_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_11(99) WHEN s_8_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_11(100) WHEN s_8_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_11(101) WHEN s_8_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_11(102) WHEN s_8_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_11(103) WHEN s_8_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_11(104) WHEN s_8_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_11(105) WHEN s_8_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_11(106) WHEN s_8_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_11(107) WHEN s_8_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_11(108) WHEN s_8_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_11(109) WHEN s_8_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_11(110) WHEN s_8_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_11(111) WHEN s_8_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_11(112) WHEN s_8_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_11(113) WHEN s_8_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_11(114) WHEN s_8_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_11(115) WHEN s_8_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_11(116) WHEN s_8_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_11(117) WHEN s_8_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_11(118) WHEN s_8_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_11(119) WHEN s_8_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_11(120) WHEN s_8_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_11(121) WHEN s_8_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_11(122) WHEN s_8_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_11(123) WHEN s_8_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_11(124) WHEN s_8_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_11(125) WHEN s_8_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_11(126) WHEN s_8_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_11(127) WHEN s_8_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_11(128) WHEN s_8_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_11(129) WHEN s_8_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_11(130) WHEN s_8_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_11(131) WHEN s_8_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_11(132) WHEN s_8_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_11(133) WHEN s_8_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_11(134) WHEN s_8_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_11(135) WHEN s_8_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_11(136) WHEN s_8_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_11(137) WHEN s_8_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_11(138) WHEN s_8_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_11(139) WHEN s_8_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_11(140) WHEN s_8_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_11(141) WHEN s_8_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_11(142) WHEN s_8_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_11(143) WHEN s_8_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_11(144) WHEN s_8_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_11(145) WHEN s_8_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_11(146) WHEN s_8_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_11(147) WHEN s_8_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_11(148) WHEN s_8_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_11(149) WHEN s_8_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_11(150) WHEN s_8_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_11(151) WHEN s_8_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_11(152) WHEN s_8_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_11(153) WHEN s_8_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_11(154) WHEN s_8_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_11(155) WHEN s_8_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_11(156) WHEN s_8_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_11(157) WHEN s_8_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_11(158) WHEN s_8_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_11(159) WHEN s_8_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_11(160) WHEN s_8_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_11(161) WHEN s_8_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_11(162) WHEN s_8_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_11(163) WHEN s_8_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_11(164) WHEN s_8_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_11(165) WHEN s_8_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_11(166) WHEN s_8_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_11(167) WHEN s_8_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_11(168) WHEN s_8_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_11(169) WHEN s_8_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_11(170) WHEN s_8_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_11(171) WHEN s_8_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_11(172) WHEN s_8_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_11(173) WHEN s_8_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_11(174) WHEN s_8_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_11(175) WHEN s_8_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_11(176) WHEN s_8_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_11(177) WHEN s_8_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_11(178) WHEN s_8_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_11(179) WHEN s_8_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_11(180) WHEN s_8_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_11(181) WHEN s_8_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_11(182) WHEN s_8_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_11(183) WHEN s_8_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_11(184) WHEN s_8_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_11(185) WHEN s_8_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_11(186) WHEN s_8_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_11(187) WHEN s_8_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_11(188) WHEN s_8_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_11(189) WHEN s_8_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_11(190) WHEN s_8_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_11(191) WHEN s_8_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_11(192) WHEN s_8_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_11(193) WHEN s_8_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_11(194) WHEN s_8_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_11(195) WHEN s_8_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_11(196) WHEN s_8_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_11(197) WHEN s_8_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_11(198) WHEN s_8_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_11(199) WHEN s_8_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_11(200) WHEN s_8_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_11(201) WHEN s_8_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_11(202) WHEN s_8_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_11(203) WHEN s_8_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_11(204) WHEN s_8_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_11(205) WHEN s_8_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_11(206) WHEN s_8_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_11(207) WHEN s_8_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_11(208) WHEN s_8_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_11(209) WHEN s_8_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_11(210) WHEN s_8_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_11(211) WHEN s_8_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_11(212) WHEN s_8_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_11(213) WHEN s_8_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_11(214) WHEN s_8_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_11(215) WHEN s_8_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_11(216) WHEN s_8_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_11(217) WHEN s_8_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_11(218) WHEN s_8_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_11(219) WHEN s_8_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_11(220) WHEN s_8_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_11(221) WHEN s_8_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_11(222) WHEN s_8_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_11(223) WHEN s_8_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_11(224) WHEN s_8_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_11(225) WHEN s_8_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_11(226) WHEN s_8_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_11(227) WHEN s_8_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_11(228) WHEN s_8_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_11(229) WHEN s_8_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_11(230) WHEN s_8_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_11(231) WHEN s_8_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_11(232) WHEN s_8_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_11(233) WHEN s_8_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_11(234) WHEN s_8_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_11(235) WHEN s_8_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_11(236) WHEN s_8_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_11(237) WHEN s_8_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_11(238) WHEN s_8_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_11(239) WHEN s_8_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_11(240) WHEN s_8_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_11(241) WHEN s_8_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_11(242) WHEN s_8_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_11(243) WHEN s_8_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_11(244) WHEN s_8_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_11(245) WHEN s_8_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_11(246) WHEN s_8_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_11(247) WHEN s_8_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_11(248) WHEN s_8_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_11(249) WHEN s_8_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_11(250) WHEN s_8_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_11(251) WHEN s_8_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_11(252) WHEN s_8_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_11(253) WHEN s_8_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_11(254) WHEN s_8_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_11(255);

  out0_145 <= out0_144 XOR s_9_1;

  b4_1 <= out0_145 XOR s_10_1;

  out0_146 <= b4_1 XOR out0_143;

  
  out0_147 <= gmul3_10(0) WHEN s_11_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_10(1) WHEN s_11_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_10(2) WHEN s_11_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_10(3) WHEN s_11_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_10(4) WHEN s_11_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_10(5) WHEN s_11_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_10(6) WHEN s_11_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_10(7) WHEN s_11_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_10(8) WHEN s_11_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_10(9) WHEN s_11_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_10(10) WHEN s_11_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_10(11) WHEN s_11_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_10(12) WHEN s_11_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_10(13) WHEN s_11_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_10(14) WHEN s_11_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_10(15) WHEN s_11_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_10(16) WHEN s_11_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_10(17) WHEN s_11_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_10(18) WHEN s_11_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_10(19) WHEN s_11_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_10(20) WHEN s_11_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_10(21) WHEN s_11_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_10(22) WHEN s_11_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_10(23) WHEN s_11_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_10(24) WHEN s_11_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_10(25) WHEN s_11_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_10(26) WHEN s_11_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_10(27) WHEN s_11_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_10(28) WHEN s_11_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_10(29) WHEN s_11_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_10(30) WHEN s_11_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_10(31) WHEN s_11_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_10(32) WHEN s_11_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_10(33) WHEN s_11_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_10(34) WHEN s_11_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_10(35) WHEN s_11_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_10(36) WHEN s_11_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_10(37) WHEN s_11_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_10(38) WHEN s_11_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_10(39) WHEN s_11_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_10(40) WHEN s_11_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_10(41) WHEN s_11_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_10(42) WHEN s_11_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_10(43) WHEN s_11_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_10(44) WHEN s_11_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_10(45) WHEN s_11_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_10(46) WHEN s_11_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_10(47) WHEN s_11_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_10(48) WHEN s_11_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_10(49) WHEN s_11_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_10(50) WHEN s_11_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_10(51) WHEN s_11_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_10(52) WHEN s_11_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_10(53) WHEN s_11_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_10(54) WHEN s_11_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_10(55) WHEN s_11_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_10(56) WHEN s_11_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_10(57) WHEN s_11_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_10(58) WHEN s_11_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_10(59) WHEN s_11_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_10(60) WHEN s_11_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_10(61) WHEN s_11_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_10(62) WHEN s_11_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_10(63) WHEN s_11_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_10(64) WHEN s_11_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_10(65) WHEN s_11_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_10(66) WHEN s_11_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_10(67) WHEN s_11_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_10(68) WHEN s_11_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_10(69) WHEN s_11_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_10(70) WHEN s_11_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_10(71) WHEN s_11_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_10(72) WHEN s_11_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_10(73) WHEN s_11_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_10(74) WHEN s_11_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_10(75) WHEN s_11_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_10(76) WHEN s_11_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_10(77) WHEN s_11_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_10(78) WHEN s_11_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_10(79) WHEN s_11_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_10(80) WHEN s_11_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_10(81) WHEN s_11_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_10(82) WHEN s_11_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_10(83) WHEN s_11_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_10(84) WHEN s_11_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_10(85) WHEN s_11_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_10(86) WHEN s_11_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_10(87) WHEN s_11_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_10(88) WHEN s_11_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_10(89) WHEN s_11_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_10(90) WHEN s_11_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_10(91) WHEN s_11_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_10(92) WHEN s_11_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_10(93) WHEN s_11_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_10(94) WHEN s_11_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_10(95) WHEN s_11_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_10(96) WHEN s_11_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_10(97) WHEN s_11_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_10(98) WHEN s_11_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_10(99) WHEN s_11_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_10(100) WHEN s_11_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_10(101) WHEN s_11_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_10(102) WHEN s_11_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_10(103) WHEN s_11_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_10(104) WHEN s_11_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_10(105) WHEN s_11_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_10(106) WHEN s_11_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_10(107) WHEN s_11_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_10(108) WHEN s_11_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_10(109) WHEN s_11_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_10(110) WHEN s_11_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_10(111) WHEN s_11_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_10(112) WHEN s_11_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_10(113) WHEN s_11_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_10(114) WHEN s_11_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_10(115) WHEN s_11_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_10(116) WHEN s_11_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_10(117) WHEN s_11_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_10(118) WHEN s_11_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_10(119) WHEN s_11_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_10(120) WHEN s_11_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_10(121) WHEN s_11_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_10(122) WHEN s_11_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_10(123) WHEN s_11_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_10(124) WHEN s_11_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_10(125) WHEN s_11_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_10(126) WHEN s_11_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_10(127) WHEN s_11_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_10(128) WHEN s_11_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_10(129) WHEN s_11_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_10(130) WHEN s_11_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_10(131) WHEN s_11_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_10(132) WHEN s_11_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_10(133) WHEN s_11_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_10(134) WHEN s_11_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_10(135) WHEN s_11_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_10(136) WHEN s_11_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_10(137) WHEN s_11_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_10(138) WHEN s_11_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_10(139) WHEN s_11_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_10(140) WHEN s_11_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_10(141) WHEN s_11_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_10(142) WHEN s_11_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_10(143) WHEN s_11_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_10(144) WHEN s_11_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_10(145) WHEN s_11_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_10(146) WHEN s_11_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_10(147) WHEN s_11_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_10(148) WHEN s_11_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_10(149) WHEN s_11_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_10(150) WHEN s_11_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_10(151) WHEN s_11_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_10(152) WHEN s_11_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_10(153) WHEN s_11_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_10(154) WHEN s_11_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_10(155) WHEN s_11_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_10(156) WHEN s_11_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_10(157) WHEN s_11_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_10(158) WHEN s_11_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_10(159) WHEN s_11_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_10(160) WHEN s_11_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_10(161) WHEN s_11_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_10(162) WHEN s_11_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_10(163) WHEN s_11_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_10(164) WHEN s_11_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_10(165) WHEN s_11_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_10(166) WHEN s_11_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_10(167) WHEN s_11_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_10(168) WHEN s_11_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_10(169) WHEN s_11_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_10(170) WHEN s_11_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_10(171) WHEN s_11_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_10(172) WHEN s_11_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_10(173) WHEN s_11_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_10(174) WHEN s_11_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_10(175) WHEN s_11_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_10(176) WHEN s_11_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_10(177) WHEN s_11_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_10(178) WHEN s_11_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_10(179) WHEN s_11_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_10(180) WHEN s_11_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_10(181) WHEN s_11_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_10(182) WHEN s_11_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_10(183) WHEN s_11_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_10(184) WHEN s_11_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_10(185) WHEN s_11_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_10(186) WHEN s_11_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_10(187) WHEN s_11_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_10(188) WHEN s_11_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_10(189) WHEN s_11_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_10(190) WHEN s_11_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_10(191) WHEN s_11_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_10(192) WHEN s_11_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_10(193) WHEN s_11_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_10(194) WHEN s_11_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_10(195) WHEN s_11_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_10(196) WHEN s_11_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_10(197) WHEN s_11_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_10(198) WHEN s_11_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_10(199) WHEN s_11_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_10(200) WHEN s_11_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_10(201) WHEN s_11_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_10(202) WHEN s_11_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_10(203) WHEN s_11_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_10(204) WHEN s_11_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_10(205) WHEN s_11_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_10(206) WHEN s_11_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_10(207) WHEN s_11_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_10(208) WHEN s_11_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_10(209) WHEN s_11_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_10(210) WHEN s_11_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_10(211) WHEN s_11_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_10(212) WHEN s_11_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_10(213) WHEN s_11_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_10(214) WHEN s_11_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_10(215) WHEN s_11_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_10(216) WHEN s_11_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_10(217) WHEN s_11_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_10(218) WHEN s_11_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_10(219) WHEN s_11_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_10(220) WHEN s_11_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_10(221) WHEN s_11_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_10(222) WHEN s_11_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_10(223) WHEN s_11_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_10(224) WHEN s_11_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_10(225) WHEN s_11_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_10(226) WHEN s_11_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_10(227) WHEN s_11_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_10(228) WHEN s_11_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_10(229) WHEN s_11_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_10(230) WHEN s_11_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_10(231) WHEN s_11_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_10(232) WHEN s_11_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_10(233) WHEN s_11_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_10(234) WHEN s_11_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_10(235) WHEN s_11_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_10(236) WHEN s_11_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_10(237) WHEN s_11_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_10(238) WHEN s_11_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_10(239) WHEN s_11_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_10(240) WHEN s_11_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_10(241) WHEN s_11_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_10(242) WHEN s_11_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_10(243) WHEN s_11_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_10(244) WHEN s_11_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_10(245) WHEN s_11_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_10(246) WHEN s_11_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_10(247) WHEN s_11_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_10(248) WHEN s_11_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_10(249) WHEN s_11_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_10(250) WHEN s_11_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_10(251) WHEN s_11_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_10(252) WHEN s_11_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_10(253) WHEN s_11_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_10(254) WHEN s_11_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_10(255);

  
  out0_148 <= gmul2_10(0) WHEN s_10_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_10(1) WHEN s_10_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_10(2) WHEN s_10_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_10(3) WHEN s_10_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_10(4) WHEN s_10_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_10(5) WHEN s_10_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_10(6) WHEN s_10_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_10(7) WHEN s_10_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_10(8) WHEN s_10_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_10(9) WHEN s_10_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_10(10) WHEN s_10_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_10(11) WHEN s_10_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_10(12) WHEN s_10_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_10(13) WHEN s_10_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_10(14) WHEN s_10_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_10(15) WHEN s_10_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_10(16) WHEN s_10_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_10(17) WHEN s_10_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_10(18) WHEN s_10_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_10(19) WHEN s_10_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_10(20) WHEN s_10_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_10(21) WHEN s_10_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_10(22) WHEN s_10_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_10(23) WHEN s_10_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_10(24) WHEN s_10_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_10(25) WHEN s_10_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_10(26) WHEN s_10_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_10(27) WHEN s_10_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_10(28) WHEN s_10_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_10(29) WHEN s_10_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_10(30) WHEN s_10_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_10(31) WHEN s_10_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_10(32) WHEN s_10_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_10(33) WHEN s_10_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_10(34) WHEN s_10_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_10(35) WHEN s_10_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_10(36) WHEN s_10_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_10(37) WHEN s_10_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_10(38) WHEN s_10_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_10(39) WHEN s_10_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_10(40) WHEN s_10_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_10(41) WHEN s_10_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_10(42) WHEN s_10_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_10(43) WHEN s_10_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_10(44) WHEN s_10_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_10(45) WHEN s_10_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_10(46) WHEN s_10_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_10(47) WHEN s_10_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_10(48) WHEN s_10_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_10(49) WHEN s_10_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_10(50) WHEN s_10_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_10(51) WHEN s_10_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_10(52) WHEN s_10_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_10(53) WHEN s_10_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_10(54) WHEN s_10_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_10(55) WHEN s_10_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_10(56) WHEN s_10_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_10(57) WHEN s_10_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_10(58) WHEN s_10_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_10(59) WHEN s_10_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_10(60) WHEN s_10_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_10(61) WHEN s_10_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_10(62) WHEN s_10_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_10(63) WHEN s_10_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_10(64) WHEN s_10_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_10(65) WHEN s_10_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_10(66) WHEN s_10_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_10(67) WHEN s_10_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_10(68) WHEN s_10_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_10(69) WHEN s_10_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_10(70) WHEN s_10_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_10(71) WHEN s_10_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_10(72) WHEN s_10_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_10(73) WHEN s_10_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_10(74) WHEN s_10_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_10(75) WHEN s_10_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_10(76) WHEN s_10_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_10(77) WHEN s_10_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_10(78) WHEN s_10_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_10(79) WHEN s_10_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_10(80) WHEN s_10_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_10(81) WHEN s_10_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_10(82) WHEN s_10_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_10(83) WHEN s_10_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_10(84) WHEN s_10_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_10(85) WHEN s_10_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_10(86) WHEN s_10_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_10(87) WHEN s_10_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_10(88) WHEN s_10_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_10(89) WHEN s_10_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_10(90) WHEN s_10_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_10(91) WHEN s_10_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_10(92) WHEN s_10_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_10(93) WHEN s_10_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_10(94) WHEN s_10_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_10(95) WHEN s_10_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_10(96) WHEN s_10_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_10(97) WHEN s_10_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_10(98) WHEN s_10_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_10(99) WHEN s_10_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_10(100) WHEN s_10_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_10(101) WHEN s_10_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_10(102) WHEN s_10_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_10(103) WHEN s_10_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_10(104) WHEN s_10_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_10(105) WHEN s_10_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_10(106) WHEN s_10_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_10(107) WHEN s_10_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_10(108) WHEN s_10_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_10(109) WHEN s_10_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_10(110) WHEN s_10_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_10(111) WHEN s_10_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_10(112) WHEN s_10_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_10(113) WHEN s_10_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_10(114) WHEN s_10_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_10(115) WHEN s_10_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_10(116) WHEN s_10_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_10(117) WHEN s_10_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_10(118) WHEN s_10_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_10(119) WHEN s_10_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_10(120) WHEN s_10_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_10(121) WHEN s_10_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_10(122) WHEN s_10_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_10(123) WHEN s_10_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_10(124) WHEN s_10_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_10(125) WHEN s_10_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_10(126) WHEN s_10_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_10(127) WHEN s_10_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_10(128) WHEN s_10_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_10(129) WHEN s_10_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_10(130) WHEN s_10_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_10(131) WHEN s_10_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_10(132) WHEN s_10_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_10(133) WHEN s_10_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_10(134) WHEN s_10_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_10(135) WHEN s_10_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_10(136) WHEN s_10_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_10(137) WHEN s_10_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_10(138) WHEN s_10_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_10(139) WHEN s_10_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_10(140) WHEN s_10_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_10(141) WHEN s_10_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_10(142) WHEN s_10_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_10(143) WHEN s_10_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_10(144) WHEN s_10_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_10(145) WHEN s_10_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_10(146) WHEN s_10_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_10(147) WHEN s_10_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_10(148) WHEN s_10_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_10(149) WHEN s_10_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_10(150) WHEN s_10_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_10(151) WHEN s_10_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_10(152) WHEN s_10_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_10(153) WHEN s_10_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_10(154) WHEN s_10_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_10(155) WHEN s_10_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_10(156) WHEN s_10_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_10(157) WHEN s_10_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_10(158) WHEN s_10_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_10(159) WHEN s_10_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_10(160) WHEN s_10_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_10(161) WHEN s_10_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_10(162) WHEN s_10_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_10(163) WHEN s_10_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_10(164) WHEN s_10_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_10(165) WHEN s_10_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_10(166) WHEN s_10_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_10(167) WHEN s_10_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_10(168) WHEN s_10_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_10(169) WHEN s_10_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_10(170) WHEN s_10_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_10(171) WHEN s_10_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_10(172) WHEN s_10_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_10(173) WHEN s_10_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_10(174) WHEN s_10_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_10(175) WHEN s_10_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_10(176) WHEN s_10_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_10(177) WHEN s_10_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_10(178) WHEN s_10_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_10(179) WHEN s_10_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_10(180) WHEN s_10_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_10(181) WHEN s_10_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_10(182) WHEN s_10_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_10(183) WHEN s_10_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_10(184) WHEN s_10_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_10(185) WHEN s_10_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_10(186) WHEN s_10_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_10(187) WHEN s_10_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_10(188) WHEN s_10_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_10(189) WHEN s_10_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_10(190) WHEN s_10_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_10(191) WHEN s_10_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_10(192) WHEN s_10_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_10(193) WHEN s_10_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_10(194) WHEN s_10_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_10(195) WHEN s_10_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_10(196) WHEN s_10_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_10(197) WHEN s_10_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_10(198) WHEN s_10_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_10(199) WHEN s_10_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_10(200) WHEN s_10_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_10(201) WHEN s_10_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_10(202) WHEN s_10_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_10(203) WHEN s_10_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_10(204) WHEN s_10_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_10(205) WHEN s_10_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_10(206) WHEN s_10_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_10(207) WHEN s_10_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_10(208) WHEN s_10_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_10(209) WHEN s_10_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_10(210) WHEN s_10_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_10(211) WHEN s_10_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_10(212) WHEN s_10_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_10(213) WHEN s_10_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_10(214) WHEN s_10_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_10(215) WHEN s_10_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_10(216) WHEN s_10_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_10(217) WHEN s_10_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_10(218) WHEN s_10_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_10(219) WHEN s_10_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_10(220) WHEN s_10_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_10(221) WHEN s_10_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_10(222) WHEN s_10_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_10(223) WHEN s_10_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_10(224) WHEN s_10_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_10(225) WHEN s_10_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_10(226) WHEN s_10_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_10(227) WHEN s_10_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_10(228) WHEN s_10_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_10(229) WHEN s_10_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_10(230) WHEN s_10_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_10(231) WHEN s_10_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_10(232) WHEN s_10_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_10(233) WHEN s_10_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_10(234) WHEN s_10_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_10(235) WHEN s_10_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_10(236) WHEN s_10_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_10(237) WHEN s_10_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_10(238) WHEN s_10_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_10(239) WHEN s_10_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_10(240) WHEN s_10_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_10(241) WHEN s_10_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_10(242) WHEN s_10_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_10(243) WHEN s_10_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_10(244) WHEN s_10_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_10(245) WHEN s_10_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_10(246) WHEN s_10_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_10(247) WHEN s_10_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_10(248) WHEN s_10_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_10(249) WHEN s_10_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_10(250) WHEN s_10_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_10(251) WHEN s_10_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_10(252) WHEN s_10_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_10(253) WHEN s_10_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_10(254) WHEN s_10_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_10(255);

  out0_149 <= s_8_1 XOR s_9_1;

  b3_1 <= out0_149 XOR out0_148;

  out0_150 <= b3_1 XOR out0_147;

  
  out0_151 <= gmul3_9(0) WHEN s_10_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_9(1) WHEN s_10_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_9(2) WHEN s_10_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_9(3) WHEN s_10_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_9(4) WHEN s_10_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_9(5) WHEN s_10_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_9(6) WHEN s_10_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_9(7) WHEN s_10_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_9(8) WHEN s_10_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_9(9) WHEN s_10_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_9(10) WHEN s_10_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_9(11) WHEN s_10_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_9(12) WHEN s_10_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_9(13) WHEN s_10_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_9(14) WHEN s_10_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_9(15) WHEN s_10_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_9(16) WHEN s_10_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_9(17) WHEN s_10_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_9(18) WHEN s_10_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_9(19) WHEN s_10_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_9(20) WHEN s_10_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_9(21) WHEN s_10_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_9(22) WHEN s_10_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_9(23) WHEN s_10_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_9(24) WHEN s_10_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_9(25) WHEN s_10_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_9(26) WHEN s_10_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_9(27) WHEN s_10_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_9(28) WHEN s_10_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_9(29) WHEN s_10_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_9(30) WHEN s_10_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_9(31) WHEN s_10_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_9(32) WHEN s_10_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_9(33) WHEN s_10_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_9(34) WHEN s_10_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_9(35) WHEN s_10_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_9(36) WHEN s_10_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_9(37) WHEN s_10_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_9(38) WHEN s_10_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_9(39) WHEN s_10_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_9(40) WHEN s_10_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_9(41) WHEN s_10_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_9(42) WHEN s_10_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_9(43) WHEN s_10_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_9(44) WHEN s_10_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_9(45) WHEN s_10_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_9(46) WHEN s_10_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_9(47) WHEN s_10_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_9(48) WHEN s_10_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_9(49) WHEN s_10_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_9(50) WHEN s_10_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_9(51) WHEN s_10_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_9(52) WHEN s_10_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_9(53) WHEN s_10_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_9(54) WHEN s_10_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_9(55) WHEN s_10_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_9(56) WHEN s_10_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_9(57) WHEN s_10_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_9(58) WHEN s_10_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_9(59) WHEN s_10_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_9(60) WHEN s_10_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_9(61) WHEN s_10_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_9(62) WHEN s_10_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_9(63) WHEN s_10_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_9(64) WHEN s_10_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_9(65) WHEN s_10_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_9(66) WHEN s_10_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_9(67) WHEN s_10_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_9(68) WHEN s_10_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_9(69) WHEN s_10_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_9(70) WHEN s_10_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_9(71) WHEN s_10_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_9(72) WHEN s_10_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_9(73) WHEN s_10_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_9(74) WHEN s_10_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_9(75) WHEN s_10_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_9(76) WHEN s_10_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_9(77) WHEN s_10_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_9(78) WHEN s_10_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_9(79) WHEN s_10_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_9(80) WHEN s_10_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_9(81) WHEN s_10_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_9(82) WHEN s_10_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_9(83) WHEN s_10_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_9(84) WHEN s_10_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_9(85) WHEN s_10_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_9(86) WHEN s_10_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_9(87) WHEN s_10_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_9(88) WHEN s_10_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_9(89) WHEN s_10_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_9(90) WHEN s_10_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_9(91) WHEN s_10_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_9(92) WHEN s_10_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_9(93) WHEN s_10_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_9(94) WHEN s_10_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_9(95) WHEN s_10_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_9(96) WHEN s_10_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_9(97) WHEN s_10_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_9(98) WHEN s_10_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_9(99) WHEN s_10_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_9(100) WHEN s_10_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_9(101) WHEN s_10_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_9(102) WHEN s_10_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_9(103) WHEN s_10_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_9(104) WHEN s_10_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_9(105) WHEN s_10_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_9(106) WHEN s_10_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_9(107) WHEN s_10_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_9(108) WHEN s_10_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_9(109) WHEN s_10_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_9(110) WHEN s_10_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_9(111) WHEN s_10_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_9(112) WHEN s_10_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_9(113) WHEN s_10_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_9(114) WHEN s_10_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_9(115) WHEN s_10_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_9(116) WHEN s_10_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_9(117) WHEN s_10_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_9(118) WHEN s_10_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_9(119) WHEN s_10_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_9(120) WHEN s_10_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_9(121) WHEN s_10_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_9(122) WHEN s_10_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_9(123) WHEN s_10_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_9(124) WHEN s_10_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_9(125) WHEN s_10_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_9(126) WHEN s_10_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_9(127) WHEN s_10_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_9(128) WHEN s_10_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_9(129) WHEN s_10_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_9(130) WHEN s_10_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_9(131) WHEN s_10_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_9(132) WHEN s_10_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_9(133) WHEN s_10_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_9(134) WHEN s_10_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_9(135) WHEN s_10_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_9(136) WHEN s_10_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_9(137) WHEN s_10_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_9(138) WHEN s_10_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_9(139) WHEN s_10_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_9(140) WHEN s_10_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_9(141) WHEN s_10_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_9(142) WHEN s_10_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_9(143) WHEN s_10_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_9(144) WHEN s_10_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_9(145) WHEN s_10_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_9(146) WHEN s_10_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_9(147) WHEN s_10_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_9(148) WHEN s_10_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_9(149) WHEN s_10_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_9(150) WHEN s_10_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_9(151) WHEN s_10_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_9(152) WHEN s_10_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_9(153) WHEN s_10_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_9(154) WHEN s_10_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_9(155) WHEN s_10_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_9(156) WHEN s_10_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_9(157) WHEN s_10_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_9(158) WHEN s_10_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_9(159) WHEN s_10_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_9(160) WHEN s_10_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_9(161) WHEN s_10_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_9(162) WHEN s_10_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_9(163) WHEN s_10_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_9(164) WHEN s_10_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_9(165) WHEN s_10_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_9(166) WHEN s_10_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_9(167) WHEN s_10_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_9(168) WHEN s_10_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_9(169) WHEN s_10_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_9(170) WHEN s_10_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_9(171) WHEN s_10_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_9(172) WHEN s_10_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_9(173) WHEN s_10_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_9(174) WHEN s_10_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_9(175) WHEN s_10_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_9(176) WHEN s_10_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_9(177) WHEN s_10_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_9(178) WHEN s_10_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_9(179) WHEN s_10_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_9(180) WHEN s_10_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_9(181) WHEN s_10_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_9(182) WHEN s_10_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_9(183) WHEN s_10_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_9(184) WHEN s_10_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_9(185) WHEN s_10_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_9(186) WHEN s_10_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_9(187) WHEN s_10_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_9(188) WHEN s_10_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_9(189) WHEN s_10_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_9(190) WHEN s_10_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_9(191) WHEN s_10_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_9(192) WHEN s_10_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_9(193) WHEN s_10_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_9(194) WHEN s_10_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_9(195) WHEN s_10_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_9(196) WHEN s_10_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_9(197) WHEN s_10_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_9(198) WHEN s_10_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_9(199) WHEN s_10_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_9(200) WHEN s_10_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_9(201) WHEN s_10_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_9(202) WHEN s_10_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_9(203) WHEN s_10_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_9(204) WHEN s_10_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_9(205) WHEN s_10_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_9(206) WHEN s_10_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_9(207) WHEN s_10_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_9(208) WHEN s_10_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_9(209) WHEN s_10_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_9(210) WHEN s_10_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_9(211) WHEN s_10_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_9(212) WHEN s_10_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_9(213) WHEN s_10_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_9(214) WHEN s_10_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_9(215) WHEN s_10_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_9(216) WHEN s_10_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_9(217) WHEN s_10_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_9(218) WHEN s_10_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_9(219) WHEN s_10_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_9(220) WHEN s_10_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_9(221) WHEN s_10_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_9(222) WHEN s_10_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_9(223) WHEN s_10_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_9(224) WHEN s_10_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_9(225) WHEN s_10_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_9(226) WHEN s_10_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_9(227) WHEN s_10_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_9(228) WHEN s_10_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_9(229) WHEN s_10_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_9(230) WHEN s_10_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_9(231) WHEN s_10_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_9(232) WHEN s_10_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_9(233) WHEN s_10_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_9(234) WHEN s_10_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_9(235) WHEN s_10_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_9(236) WHEN s_10_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_9(237) WHEN s_10_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_9(238) WHEN s_10_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_9(239) WHEN s_10_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_9(240) WHEN s_10_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_9(241) WHEN s_10_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_9(242) WHEN s_10_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_9(243) WHEN s_10_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_9(244) WHEN s_10_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_9(245) WHEN s_10_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_9(246) WHEN s_10_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_9(247) WHEN s_10_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_9(248) WHEN s_10_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_9(249) WHEN s_10_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_9(250) WHEN s_10_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_9(251) WHEN s_10_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_9(252) WHEN s_10_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_9(253) WHEN s_10_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_9(254) WHEN s_10_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_9(255);

  
  out0_152 <= gmul2_9(0) WHEN s_9_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_9(1) WHEN s_9_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_9(2) WHEN s_9_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_9(3) WHEN s_9_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_9(4) WHEN s_9_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_9(5) WHEN s_9_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_9(6) WHEN s_9_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_9(7) WHEN s_9_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_9(8) WHEN s_9_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_9(9) WHEN s_9_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_9(10) WHEN s_9_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_9(11) WHEN s_9_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_9(12) WHEN s_9_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_9(13) WHEN s_9_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_9(14) WHEN s_9_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_9(15) WHEN s_9_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_9(16) WHEN s_9_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_9(17) WHEN s_9_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_9(18) WHEN s_9_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_9(19) WHEN s_9_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_9(20) WHEN s_9_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_9(21) WHEN s_9_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_9(22) WHEN s_9_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_9(23) WHEN s_9_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_9(24) WHEN s_9_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_9(25) WHEN s_9_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_9(26) WHEN s_9_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_9(27) WHEN s_9_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_9(28) WHEN s_9_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_9(29) WHEN s_9_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_9(30) WHEN s_9_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_9(31) WHEN s_9_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_9(32) WHEN s_9_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_9(33) WHEN s_9_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_9(34) WHEN s_9_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_9(35) WHEN s_9_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_9(36) WHEN s_9_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_9(37) WHEN s_9_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_9(38) WHEN s_9_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_9(39) WHEN s_9_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_9(40) WHEN s_9_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_9(41) WHEN s_9_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_9(42) WHEN s_9_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_9(43) WHEN s_9_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_9(44) WHEN s_9_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_9(45) WHEN s_9_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_9(46) WHEN s_9_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_9(47) WHEN s_9_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_9(48) WHEN s_9_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_9(49) WHEN s_9_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_9(50) WHEN s_9_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_9(51) WHEN s_9_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_9(52) WHEN s_9_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_9(53) WHEN s_9_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_9(54) WHEN s_9_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_9(55) WHEN s_9_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_9(56) WHEN s_9_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_9(57) WHEN s_9_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_9(58) WHEN s_9_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_9(59) WHEN s_9_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_9(60) WHEN s_9_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_9(61) WHEN s_9_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_9(62) WHEN s_9_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_9(63) WHEN s_9_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_9(64) WHEN s_9_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_9(65) WHEN s_9_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_9(66) WHEN s_9_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_9(67) WHEN s_9_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_9(68) WHEN s_9_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_9(69) WHEN s_9_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_9(70) WHEN s_9_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_9(71) WHEN s_9_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_9(72) WHEN s_9_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_9(73) WHEN s_9_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_9(74) WHEN s_9_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_9(75) WHEN s_9_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_9(76) WHEN s_9_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_9(77) WHEN s_9_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_9(78) WHEN s_9_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_9(79) WHEN s_9_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_9(80) WHEN s_9_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_9(81) WHEN s_9_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_9(82) WHEN s_9_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_9(83) WHEN s_9_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_9(84) WHEN s_9_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_9(85) WHEN s_9_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_9(86) WHEN s_9_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_9(87) WHEN s_9_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_9(88) WHEN s_9_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_9(89) WHEN s_9_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_9(90) WHEN s_9_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_9(91) WHEN s_9_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_9(92) WHEN s_9_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_9(93) WHEN s_9_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_9(94) WHEN s_9_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_9(95) WHEN s_9_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_9(96) WHEN s_9_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_9(97) WHEN s_9_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_9(98) WHEN s_9_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_9(99) WHEN s_9_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_9(100) WHEN s_9_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_9(101) WHEN s_9_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_9(102) WHEN s_9_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_9(103) WHEN s_9_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_9(104) WHEN s_9_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_9(105) WHEN s_9_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_9(106) WHEN s_9_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_9(107) WHEN s_9_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_9(108) WHEN s_9_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_9(109) WHEN s_9_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_9(110) WHEN s_9_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_9(111) WHEN s_9_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_9(112) WHEN s_9_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_9(113) WHEN s_9_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_9(114) WHEN s_9_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_9(115) WHEN s_9_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_9(116) WHEN s_9_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_9(117) WHEN s_9_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_9(118) WHEN s_9_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_9(119) WHEN s_9_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_9(120) WHEN s_9_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_9(121) WHEN s_9_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_9(122) WHEN s_9_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_9(123) WHEN s_9_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_9(124) WHEN s_9_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_9(125) WHEN s_9_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_9(126) WHEN s_9_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_9(127) WHEN s_9_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_9(128) WHEN s_9_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_9(129) WHEN s_9_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_9(130) WHEN s_9_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_9(131) WHEN s_9_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_9(132) WHEN s_9_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_9(133) WHEN s_9_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_9(134) WHEN s_9_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_9(135) WHEN s_9_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_9(136) WHEN s_9_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_9(137) WHEN s_9_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_9(138) WHEN s_9_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_9(139) WHEN s_9_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_9(140) WHEN s_9_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_9(141) WHEN s_9_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_9(142) WHEN s_9_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_9(143) WHEN s_9_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_9(144) WHEN s_9_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_9(145) WHEN s_9_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_9(146) WHEN s_9_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_9(147) WHEN s_9_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_9(148) WHEN s_9_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_9(149) WHEN s_9_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_9(150) WHEN s_9_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_9(151) WHEN s_9_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_9(152) WHEN s_9_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_9(153) WHEN s_9_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_9(154) WHEN s_9_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_9(155) WHEN s_9_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_9(156) WHEN s_9_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_9(157) WHEN s_9_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_9(158) WHEN s_9_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_9(159) WHEN s_9_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_9(160) WHEN s_9_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_9(161) WHEN s_9_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_9(162) WHEN s_9_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_9(163) WHEN s_9_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_9(164) WHEN s_9_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_9(165) WHEN s_9_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_9(166) WHEN s_9_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_9(167) WHEN s_9_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_9(168) WHEN s_9_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_9(169) WHEN s_9_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_9(170) WHEN s_9_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_9(171) WHEN s_9_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_9(172) WHEN s_9_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_9(173) WHEN s_9_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_9(174) WHEN s_9_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_9(175) WHEN s_9_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_9(176) WHEN s_9_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_9(177) WHEN s_9_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_9(178) WHEN s_9_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_9(179) WHEN s_9_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_9(180) WHEN s_9_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_9(181) WHEN s_9_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_9(182) WHEN s_9_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_9(183) WHEN s_9_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_9(184) WHEN s_9_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_9(185) WHEN s_9_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_9(186) WHEN s_9_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_9(187) WHEN s_9_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_9(188) WHEN s_9_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_9(189) WHEN s_9_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_9(190) WHEN s_9_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_9(191) WHEN s_9_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_9(192) WHEN s_9_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_9(193) WHEN s_9_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_9(194) WHEN s_9_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_9(195) WHEN s_9_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_9(196) WHEN s_9_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_9(197) WHEN s_9_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_9(198) WHEN s_9_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_9(199) WHEN s_9_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_9(200) WHEN s_9_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_9(201) WHEN s_9_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_9(202) WHEN s_9_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_9(203) WHEN s_9_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_9(204) WHEN s_9_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_9(205) WHEN s_9_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_9(206) WHEN s_9_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_9(207) WHEN s_9_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_9(208) WHEN s_9_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_9(209) WHEN s_9_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_9(210) WHEN s_9_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_9(211) WHEN s_9_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_9(212) WHEN s_9_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_9(213) WHEN s_9_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_9(214) WHEN s_9_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_9(215) WHEN s_9_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_9(216) WHEN s_9_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_9(217) WHEN s_9_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_9(218) WHEN s_9_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_9(219) WHEN s_9_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_9(220) WHEN s_9_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_9(221) WHEN s_9_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_9(222) WHEN s_9_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_9(223) WHEN s_9_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_9(224) WHEN s_9_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_9(225) WHEN s_9_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_9(226) WHEN s_9_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_9(227) WHEN s_9_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_9(228) WHEN s_9_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_9(229) WHEN s_9_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_9(230) WHEN s_9_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_9(231) WHEN s_9_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_9(232) WHEN s_9_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_9(233) WHEN s_9_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_9(234) WHEN s_9_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_9(235) WHEN s_9_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_9(236) WHEN s_9_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_9(237) WHEN s_9_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_9(238) WHEN s_9_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_9(239) WHEN s_9_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_9(240) WHEN s_9_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_9(241) WHEN s_9_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_9(242) WHEN s_9_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_9(243) WHEN s_9_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_9(244) WHEN s_9_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_9(245) WHEN s_9_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_9(246) WHEN s_9_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_9(247) WHEN s_9_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_9(248) WHEN s_9_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_9(249) WHEN s_9_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_9(250) WHEN s_9_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_9(251) WHEN s_9_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_9(252) WHEN s_9_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_9(253) WHEN s_9_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_9(254) WHEN s_9_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_9(255);

  out0_153 <= s_8_1 XOR out0_152;

  b2_1 <= out0_153 XOR out0_151;

  out0_154 <= b2_1 XOR s_11_1;

  s_11_1 <= s_s_5(11);

  s_10_1 <= s_s_5(10);

  s_9_1 <= s_s_5(9);

  
  out0_155 <= gmul3_8(0) WHEN s_9_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_8(1) WHEN s_9_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_8(2) WHEN s_9_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_8(3) WHEN s_9_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_8(4) WHEN s_9_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_8(5) WHEN s_9_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_8(6) WHEN s_9_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_8(7) WHEN s_9_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_8(8) WHEN s_9_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_8(9) WHEN s_9_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_8(10) WHEN s_9_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_8(11) WHEN s_9_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_8(12) WHEN s_9_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_8(13) WHEN s_9_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_8(14) WHEN s_9_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_8(15) WHEN s_9_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_8(16) WHEN s_9_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_8(17) WHEN s_9_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_8(18) WHEN s_9_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_8(19) WHEN s_9_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_8(20) WHEN s_9_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_8(21) WHEN s_9_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_8(22) WHEN s_9_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_8(23) WHEN s_9_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_8(24) WHEN s_9_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_8(25) WHEN s_9_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_8(26) WHEN s_9_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_8(27) WHEN s_9_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_8(28) WHEN s_9_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_8(29) WHEN s_9_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_8(30) WHEN s_9_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_8(31) WHEN s_9_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_8(32) WHEN s_9_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_8(33) WHEN s_9_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_8(34) WHEN s_9_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_8(35) WHEN s_9_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_8(36) WHEN s_9_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_8(37) WHEN s_9_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_8(38) WHEN s_9_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_8(39) WHEN s_9_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_8(40) WHEN s_9_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_8(41) WHEN s_9_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_8(42) WHEN s_9_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_8(43) WHEN s_9_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_8(44) WHEN s_9_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_8(45) WHEN s_9_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_8(46) WHEN s_9_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_8(47) WHEN s_9_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_8(48) WHEN s_9_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_8(49) WHEN s_9_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_8(50) WHEN s_9_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_8(51) WHEN s_9_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_8(52) WHEN s_9_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_8(53) WHEN s_9_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_8(54) WHEN s_9_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_8(55) WHEN s_9_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_8(56) WHEN s_9_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_8(57) WHEN s_9_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_8(58) WHEN s_9_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_8(59) WHEN s_9_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_8(60) WHEN s_9_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_8(61) WHEN s_9_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_8(62) WHEN s_9_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_8(63) WHEN s_9_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_8(64) WHEN s_9_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_8(65) WHEN s_9_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_8(66) WHEN s_9_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_8(67) WHEN s_9_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_8(68) WHEN s_9_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_8(69) WHEN s_9_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_8(70) WHEN s_9_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_8(71) WHEN s_9_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_8(72) WHEN s_9_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_8(73) WHEN s_9_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_8(74) WHEN s_9_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_8(75) WHEN s_9_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_8(76) WHEN s_9_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_8(77) WHEN s_9_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_8(78) WHEN s_9_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_8(79) WHEN s_9_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_8(80) WHEN s_9_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_8(81) WHEN s_9_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_8(82) WHEN s_9_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_8(83) WHEN s_9_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_8(84) WHEN s_9_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_8(85) WHEN s_9_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_8(86) WHEN s_9_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_8(87) WHEN s_9_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_8(88) WHEN s_9_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_8(89) WHEN s_9_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_8(90) WHEN s_9_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_8(91) WHEN s_9_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_8(92) WHEN s_9_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_8(93) WHEN s_9_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_8(94) WHEN s_9_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_8(95) WHEN s_9_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_8(96) WHEN s_9_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_8(97) WHEN s_9_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_8(98) WHEN s_9_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_8(99) WHEN s_9_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_8(100) WHEN s_9_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_8(101) WHEN s_9_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_8(102) WHEN s_9_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_8(103) WHEN s_9_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_8(104) WHEN s_9_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_8(105) WHEN s_9_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_8(106) WHEN s_9_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_8(107) WHEN s_9_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_8(108) WHEN s_9_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_8(109) WHEN s_9_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_8(110) WHEN s_9_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_8(111) WHEN s_9_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_8(112) WHEN s_9_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_8(113) WHEN s_9_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_8(114) WHEN s_9_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_8(115) WHEN s_9_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_8(116) WHEN s_9_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_8(117) WHEN s_9_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_8(118) WHEN s_9_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_8(119) WHEN s_9_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_8(120) WHEN s_9_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_8(121) WHEN s_9_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_8(122) WHEN s_9_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_8(123) WHEN s_9_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_8(124) WHEN s_9_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_8(125) WHEN s_9_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_8(126) WHEN s_9_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_8(127) WHEN s_9_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_8(128) WHEN s_9_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_8(129) WHEN s_9_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_8(130) WHEN s_9_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_8(131) WHEN s_9_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_8(132) WHEN s_9_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_8(133) WHEN s_9_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_8(134) WHEN s_9_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_8(135) WHEN s_9_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_8(136) WHEN s_9_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_8(137) WHEN s_9_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_8(138) WHEN s_9_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_8(139) WHEN s_9_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_8(140) WHEN s_9_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_8(141) WHEN s_9_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_8(142) WHEN s_9_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_8(143) WHEN s_9_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_8(144) WHEN s_9_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_8(145) WHEN s_9_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_8(146) WHEN s_9_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_8(147) WHEN s_9_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_8(148) WHEN s_9_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_8(149) WHEN s_9_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_8(150) WHEN s_9_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_8(151) WHEN s_9_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_8(152) WHEN s_9_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_8(153) WHEN s_9_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_8(154) WHEN s_9_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_8(155) WHEN s_9_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_8(156) WHEN s_9_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_8(157) WHEN s_9_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_8(158) WHEN s_9_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_8(159) WHEN s_9_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_8(160) WHEN s_9_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_8(161) WHEN s_9_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_8(162) WHEN s_9_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_8(163) WHEN s_9_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_8(164) WHEN s_9_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_8(165) WHEN s_9_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_8(166) WHEN s_9_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_8(167) WHEN s_9_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_8(168) WHEN s_9_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_8(169) WHEN s_9_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_8(170) WHEN s_9_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_8(171) WHEN s_9_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_8(172) WHEN s_9_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_8(173) WHEN s_9_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_8(174) WHEN s_9_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_8(175) WHEN s_9_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_8(176) WHEN s_9_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_8(177) WHEN s_9_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_8(178) WHEN s_9_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_8(179) WHEN s_9_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_8(180) WHEN s_9_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_8(181) WHEN s_9_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_8(182) WHEN s_9_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_8(183) WHEN s_9_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_8(184) WHEN s_9_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_8(185) WHEN s_9_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_8(186) WHEN s_9_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_8(187) WHEN s_9_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_8(188) WHEN s_9_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_8(189) WHEN s_9_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_8(190) WHEN s_9_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_8(191) WHEN s_9_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_8(192) WHEN s_9_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_8(193) WHEN s_9_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_8(194) WHEN s_9_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_8(195) WHEN s_9_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_8(196) WHEN s_9_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_8(197) WHEN s_9_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_8(198) WHEN s_9_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_8(199) WHEN s_9_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_8(200) WHEN s_9_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_8(201) WHEN s_9_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_8(202) WHEN s_9_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_8(203) WHEN s_9_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_8(204) WHEN s_9_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_8(205) WHEN s_9_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_8(206) WHEN s_9_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_8(207) WHEN s_9_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_8(208) WHEN s_9_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_8(209) WHEN s_9_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_8(210) WHEN s_9_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_8(211) WHEN s_9_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_8(212) WHEN s_9_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_8(213) WHEN s_9_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_8(214) WHEN s_9_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_8(215) WHEN s_9_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_8(216) WHEN s_9_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_8(217) WHEN s_9_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_8(218) WHEN s_9_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_8(219) WHEN s_9_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_8(220) WHEN s_9_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_8(221) WHEN s_9_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_8(222) WHEN s_9_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_8(223) WHEN s_9_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_8(224) WHEN s_9_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_8(225) WHEN s_9_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_8(226) WHEN s_9_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_8(227) WHEN s_9_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_8(228) WHEN s_9_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_8(229) WHEN s_9_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_8(230) WHEN s_9_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_8(231) WHEN s_9_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_8(232) WHEN s_9_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_8(233) WHEN s_9_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_8(234) WHEN s_9_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_8(235) WHEN s_9_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_8(236) WHEN s_9_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_8(237) WHEN s_9_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_8(238) WHEN s_9_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_8(239) WHEN s_9_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_8(240) WHEN s_9_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_8(241) WHEN s_9_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_8(242) WHEN s_9_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_8(243) WHEN s_9_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_8(244) WHEN s_9_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_8(245) WHEN s_9_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_8(246) WHEN s_9_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_8(247) WHEN s_9_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_8(248) WHEN s_9_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_8(249) WHEN s_9_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_8(250) WHEN s_9_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_8(251) WHEN s_9_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_8(252) WHEN s_9_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_8(253) WHEN s_9_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_8(254) WHEN s_9_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_8(255);

  s_8_1 <= s_s_5(8);

  
  out0_156 <= gmul2_8(0) WHEN s_8_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_8(1) WHEN s_8_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_8(2) WHEN s_8_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_8(3) WHEN s_8_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_8(4) WHEN s_8_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_8(5) WHEN s_8_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_8(6) WHEN s_8_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_8(7) WHEN s_8_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_8(8) WHEN s_8_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_8(9) WHEN s_8_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_8(10) WHEN s_8_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_8(11) WHEN s_8_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_8(12) WHEN s_8_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_8(13) WHEN s_8_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_8(14) WHEN s_8_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_8(15) WHEN s_8_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_8(16) WHEN s_8_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_8(17) WHEN s_8_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_8(18) WHEN s_8_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_8(19) WHEN s_8_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_8(20) WHEN s_8_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_8(21) WHEN s_8_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_8(22) WHEN s_8_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_8(23) WHEN s_8_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_8(24) WHEN s_8_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_8(25) WHEN s_8_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_8(26) WHEN s_8_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_8(27) WHEN s_8_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_8(28) WHEN s_8_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_8(29) WHEN s_8_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_8(30) WHEN s_8_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_8(31) WHEN s_8_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_8(32) WHEN s_8_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_8(33) WHEN s_8_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_8(34) WHEN s_8_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_8(35) WHEN s_8_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_8(36) WHEN s_8_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_8(37) WHEN s_8_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_8(38) WHEN s_8_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_8(39) WHEN s_8_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_8(40) WHEN s_8_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_8(41) WHEN s_8_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_8(42) WHEN s_8_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_8(43) WHEN s_8_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_8(44) WHEN s_8_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_8(45) WHEN s_8_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_8(46) WHEN s_8_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_8(47) WHEN s_8_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_8(48) WHEN s_8_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_8(49) WHEN s_8_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_8(50) WHEN s_8_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_8(51) WHEN s_8_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_8(52) WHEN s_8_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_8(53) WHEN s_8_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_8(54) WHEN s_8_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_8(55) WHEN s_8_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_8(56) WHEN s_8_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_8(57) WHEN s_8_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_8(58) WHEN s_8_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_8(59) WHEN s_8_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_8(60) WHEN s_8_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_8(61) WHEN s_8_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_8(62) WHEN s_8_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_8(63) WHEN s_8_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_8(64) WHEN s_8_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_8(65) WHEN s_8_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_8(66) WHEN s_8_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_8(67) WHEN s_8_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_8(68) WHEN s_8_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_8(69) WHEN s_8_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_8(70) WHEN s_8_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_8(71) WHEN s_8_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_8(72) WHEN s_8_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_8(73) WHEN s_8_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_8(74) WHEN s_8_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_8(75) WHEN s_8_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_8(76) WHEN s_8_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_8(77) WHEN s_8_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_8(78) WHEN s_8_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_8(79) WHEN s_8_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_8(80) WHEN s_8_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_8(81) WHEN s_8_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_8(82) WHEN s_8_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_8(83) WHEN s_8_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_8(84) WHEN s_8_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_8(85) WHEN s_8_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_8(86) WHEN s_8_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_8(87) WHEN s_8_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_8(88) WHEN s_8_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_8(89) WHEN s_8_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_8(90) WHEN s_8_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_8(91) WHEN s_8_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_8(92) WHEN s_8_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_8(93) WHEN s_8_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_8(94) WHEN s_8_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_8(95) WHEN s_8_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_8(96) WHEN s_8_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_8(97) WHEN s_8_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_8(98) WHEN s_8_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_8(99) WHEN s_8_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_8(100) WHEN s_8_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_8(101) WHEN s_8_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_8(102) WHEN s_8_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_8(103) WHEN s_8_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_8(104) WHEN s_8_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_8(105) WHEN s_8_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_8(106) WHEN s_8_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_8(107) WHEN s_8_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_8(108) WHEN s_8_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_8(109) WHEN s_8_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_8(110) WHEN s_8_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_8(111) WHEN s_8_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_8(112) WHEN s_8_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_8(113) WHEN s_8_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_8(114) WHEN s_8_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_8(115) WHEN s_8_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_8(116) WHEN s_8_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_8(117) WHEN s_8_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_8(118) WHEN s_8_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_8(119) WHEN s_8_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_8(120) WHEN s_8_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_8(121) WHEN s_8_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_8(122) WHEN s_8_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_8(123) WHEN s_8_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_8(124) WHEN s_8_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_8(125) WHEN s_8_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_8(126) WHEN s_8_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_8(127) WHEN s_8_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_8(128) WHEN s_8_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_8(129) WHEN s_8_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_8(130) WHEN s_8_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_8(131) WHEN s_8_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_8(132) WHEN s_8_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_8(133) WHEN s_8_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_8(134) WHEN s_8_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_8(135) WHEN s_8_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_8(136) WHEN s_8_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_8(137) WHEN s_8_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_8(138) WHEN s_8_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_8(139) WHEN s_8_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_8(140) WHEN s_8_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_8(141) WHEN s_8_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_8(142) WHEN s_8_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_8(143) WHEN s_8_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_8(144) WHEN s_8_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_8(145) WHEN s_8_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_8(146) WHEN s_8_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_8(147) WHEN s_8_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_8(148) WHEN s_8_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_8(149) WHEN s_8_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_8(150) WHEN s_8_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_8(151) WHEN s_8_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_8(152) WHEN s_8_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_8(153) WHEN s_8_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_8(154) WHEN s_8_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_8(155) WHEN s_8_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_8(156) WHEN s_8_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_8(157) WHEN s_8_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_8(158) WHEN s_8_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_8(159) WHEN s_8_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_8(160) WHEN s_8_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_8(161) WHEN s_8_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_8(162) WHEN s_8_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_8(163) WHEN s_8_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_8(164) WHEN s_8_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_8(165) WHEN s_8_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_8(166) WHEN s_8_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_8(167) WHEN s_8_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_8(168) WHEN s_8_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_8(169) WHEN s_8_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_8(170) WHEN s_8_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_8(171) WHEN s_8_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_8(172) WHEN s_8_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_8(173) WHEN s_8_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_8(174) WHEN s_8_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_8(175) WHEN s_8_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_8(176) WHEN s_8_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_8(177) WHEN s_8_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_8(178) WHEN s_8_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_8(179) WHEN s_8_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_8(180) WHEN s_8_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_8(181) WHEN s_8_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_8(182) WHEN s_8_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_8(183) WHEN s_8_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_8(184) WHEN s_8_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_8(185) WHEN s_8_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_8(186) WHEN s_8_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_8(187) WHEN s_8_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_8(188) WHEN s_8_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_8(189) WHEN s_8_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_8(190) WHEN s_8_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_8(191) WHEN s_8_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_8(192) WHEN s_8_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_8(193) WHEN s_8_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_8(194) WHEN s_8_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_8(195) WHEN s_8_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_8(196) WHEN s_8_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_8(197) WHEN s_8_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_8(198) WHEN s_8_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_8(199) WHEN s_8_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_8(200) WHEN s_8_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_8(201) WHEN s_8_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_8(202) WHEN s_8_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_8(203) WHEN s_8_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_8(204) WHEN s_8_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_8(205) WHEN s_8_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_8(206) WHEN s_8_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_8(207) WHEN s_8_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_8(208) WHEN s_8_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_8(209) WHEN s_8_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_8(210) WHEN s_8_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_8(211) WHEN s_8_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_8(212) WHEN s_8_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_8(213) WHEN s_8_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_8(214) WHEN s_8_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_8(215) WHEN s_8_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_8(216) WHEN s_8_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_8(217) WHEN s_8_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_8(218) WHEN s_8_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_8(219) WHEN s_8_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_8(220) WHEN s_8_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_8(221) WHEN s_8_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_8(222) WHEN s_8_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_8(223) WHEN s_8_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_8(224) WHEN s_8_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_8(225) WHEN s_8_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_8(226) WHEN s_8_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_8(227) WHEN s_8_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_8(228) WHEN s_8_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_8(229) WHEN s_8_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_8(230) WHEN s_8_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_8(231) WHEN s_8_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_8(232) WHEN s_8_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_8(233) WHEN s_8_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_8(234) WHEN s_8_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_8(235) WHEN s_8_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_8(236) WHEN s_8_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_8(237) WHEN s_8_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_8(238) WHEN s_8_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_8(239) WHEN s_8_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_8(240) WHEN s_8_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_8(241) WHEN s_8_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_8(242) WHEN s_8_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_8(243) WHEN s_8_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_8(244) WHEN s_8_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_8(245) WHEN s_8_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_8(246) WHEN s_8_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_8(247) WHEN s_8_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_8(248) WHEN s_8_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_8(249) WHEN s_8_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_8(250) WHEN s_8_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_8(251) WHEN s_8_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_8(252) WHEN s_8_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_8(253) WHEN s_8_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_8(254) WHEN s_8_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_8(255);

  out0_157 <= out0_156 XOR out0_155;

  b1_1 <= out0_157 XOR s_10_1;

  out0_158 <= b1_1 XOR s_11_1;

  
  out0_159 <= gmul2_7(0) WHEN s_7_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_7(1) WHEN s_7_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_7(2) WHEN s_7_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_7(3) WHEN s_7_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_7(4) WHEN s_7_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_7(5) WHEN s_7_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_7(6) WHEN s_7_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_7(7) WHEN s_7_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_7(8) WHEN s_7_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_7(9) WHEN s_7_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_7(10) WHEN s_7_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_7(11) WHEN s_7_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_7(12) WHEN s_7_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_7(13) WHEN s_7_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_7(14) WHEN s_7_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_7(15) WHEN s_7_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_7(16) WHEN s_7_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_7(17) WHEN s_7_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_7(18) WHEN s_7_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_7(19) WHEN s_7_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_7(20) WHEN s_7_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_7(21) WHEN s_7_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_7(22) WHEN s_7_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_7(23) WHEN s_7_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_7(24) WHEN s_7_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_7(25) WHEN s_7_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_7(26) WHEN s_7_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_7(27) WHEN s_7_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_7(28) WHEN s_7_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_7(29) WHEN s_7_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_7(30) WHEN s_7_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_7(31) WHEN s_7_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_7(32) WHEN s_7_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_7(33) WHEN s_7_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_7(34) WHEN s_7_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_7(35) WHEN s_7_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_7(36) WHEN s_7_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_7(37) WHEN s_7_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_7(38) WHEN s_7_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_7(39) WHEN s_7_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_7(40) WHEN s_7_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_7(41) WHEN s_7_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_7(42) WHEN s_7_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_7(43) WHEN s_7_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_7(44) WHEN s_7_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_7(45) WHEN s_7_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_7(46) WHEN s_7_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_7(47) WHEN s_7_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_7(48) WHEN s_7_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_7(49) WHEN s_7_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_7(50) WHEN s_7_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_7(51) WHEN s_7_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_7(52) WHEN s_7_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_7(53) WHEN s_7_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_7(54) WHEN s_7_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_7(55) WHEN s_7_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_7(56) WHEN s_7_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_7(57) WHEN s_7_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_7(58) WHEN s_7_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_7(59) WHEN s_7_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_7(60) WHEN s_7_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_7(61) WHEN s_7_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_7(62) WHEN s_7_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_7(63) WHEN s_7_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_7(64) WHEN s_7_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_7(65) WHEN s_7_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_7(66) WHEN s_7_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_7(67) WHEN s_7_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_7(68) WHEN s_7_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_7(69) WHEN s_7_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_7(70) WHEN s_7_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_7(71) WHEN s_7_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_7(72) WHEN s_7_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_7(73) WHEN s_7_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_7(74) WHEN s_7_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_7(75) WHEN s_7_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_7(76) WHEN s_7_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_7(77) WHEN s_7_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_7(78) WHEN s_7_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_7(79) WHEN s_7_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_7(80) WHEN s_7_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_7(81) WHEN s_7_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_7(82) WHEN s_7_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_7(83) WHEN s_7_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_7(84) WHEN s_7_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_7(85) WHEN s_7_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_7(86) WHEN s_7_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_7(87) WHEN s_7_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_7(88) WHEN s_7_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_7(89) WHEN s_7_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_7(90) WHEN s_7_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_7(91) WHEN s_7_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_7(92) WHEN s_7_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_7(93) WHEN s_7_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_7(94) WHEN s_7_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_7(95) WHEN s_7_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_7(96) WHEN s_7_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_7(97) WHEN s_7_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_7(98) WHEN s_7_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_7(99) WHEN s_7_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_7(100) WHEN s_7_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_7(101) WHEN s_7_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_7(102) WHEN s_7_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_7(103) WHEN s_7_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_7(104) WHEN s_7_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_7(105) WHEN s_7_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_7(106) WHEN s_7_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_7(107) WHEN s_7_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_7(108) WHEN s_7_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_7(109) WHEN s_7_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_7(110) WHEN s_7_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_7(111) WHEN s_7_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_7(112) WHEN s_7_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_7(113) WHEN s_7_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_7(114) WHEN s_7_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_7(115) WHEN s_7_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_7(116) WHEN s_7_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_7(117) WHEN s_7_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_7(118) WHEN s_7_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_7(119) WHEN s_7_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_7(120) WHEN s_7_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_7(121) WHEN s_7_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_7(122) WHEN s_7_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_7(123) WHEN s_7_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_7(124) WHEN s_7_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_7(125) WHEN s_7_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_7(126) WHEN s_7_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_7(127) WHEN s_7_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_7(128) WHEN s_7_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_7(129) WHEN s_7_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_7(130) WHEN s_7_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_7(131) WHEN s_7_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_7(132) WHEN s_7_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_7(133) WHEN s_7_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_7(134) WHEN s_7_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_7(135) WHEN s_7_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_7(136) WHEN s_7_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_7(137) WHEN s_7_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_7(138) WHEN s_7_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_7(139) WHEN s_7_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_7(140) WHEN s_7_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_7(141) WHEN s_7_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_7(142) WHEN s_7_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_7(143) WHEN s_7_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_7(144) WHEN s_7_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_7(145) WHEN s_7_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_7(146) WHEN s_7_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_7(147) WHEN s_7_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_7(148) WHEN s_7_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_7(149) WHEN s_7_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_7(150) WHEN s_7_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_7(151) WHEN s_7_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_7(152) WHEN s_7_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_7(153) WHEN s_7_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_7(154) WHEN s_7_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_7(155) WHEN s_7_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_7(156) WHEN s_7_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_7(157) WHEN s_7_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_7(158) WHEN s_7_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_7(159) WHEN s_7_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_7(160) WHEN s_7_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_7(161) WHEN s_7_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_7(162) WHEN s_7_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_7(163) WHEN s_7_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_7(164) WHEN s_7_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_7(165) WHEN s_7_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_7(166) WHEN s_7_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_7(167) WHEN s_7_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_7(168) WHEN s_7_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_7(169) WHEN s_7_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_7(170) WHEN s_7_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_7(171) WHEN s_7_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_7(172) WHEN s_7_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_7(173) WHEN s_7_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_7(174) WHEN s_7_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_7(175) WHEN s_7_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_7(176) WHEN s_7_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_7(177) WHEN s_7_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_7(178) WHEN s_7_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_7(179) WHEN s_7_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_7(180) WHEN s_7_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_7(181) WHEN s_7_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_7(182) WHEN s_7_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_7(183) WHEN s_7_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_7(184) WHEN s_7_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_7(185) WHEN s_7_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_7(186) WHEN s_7_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_7(187) WHEN s_7_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_7(188) WHEN s_7_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_7(189) WHEN s_7_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_7(190) WHEN s_7_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_7(191) WHEN s_7_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_7(192) WHEN s_7_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_7(193) WHEN s_7_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_7(194) WHEN s_7_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_7(195) WHEN s_7_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_7(196) WHEN s_7_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_7(197) WHEN s_7_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_7(198) WHEN s_7_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_7(199) WHEN s_7_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_7(200) WHEN s_7_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_7(201) WHEN s_7_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_7(202) WHEN s_7_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_7(203) WHEN s_7_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_7(204) WHEN s_7_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_7(205) WHEN s_7_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_7(206) WHEN s_7_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_7(207) WHEN s_7_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_7(208) WHEN s_7_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_7(209) WHEN s_7_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_7(210) WHEN s_7_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_7(211) WHEN s_7_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_7(212) WHEN s_7_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_7(213) WHEN s_7_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_7(214) WHEN s_7_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_7(215) WHEN s_7_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_7(216) WHEN s_7_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_7(217) WHEN s_7_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_7(218) WHEN s_7_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_7(219) WHEN s_7_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_7(220) WHEN s_7_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_7(221) WHEN s_7_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_7(222) WHEN s_7_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_7(223) WHEN s_7_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_7(224) WHEN s_7_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_7(225) WHEN s_7_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_7(226) WHEN s_7_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_7(227) WHEN s_7_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_7(228) WHEN s_7_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_7(229) WHEN s_7_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_7(230) WHEN s_7_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_7(231) WHEN s_7_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_7(232) WHEN s_7_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_7(233) WHEN s_7_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_7(234) WHEN s_7_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_7(235) WHEN s_7_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_7(236) WHEN s_7_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_7(237) WHEN s_7_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_7(238) WHEN s_7_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_7(239) WHEN s_7_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_7(240) WHEN s_7_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_7(241) WHEN s_7_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_7(242) WHEN s_7_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_7(243) WHEN s_7_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_7(244) WHEN s_7_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_7(245) WHEN s_7_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_7(246) WHEN s_7_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_7(247) WHEN s_7_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_7(248) WHEN s_7_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_7(249) WHEN s_7_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_7(250) WHEN s_7_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_7(251) WHEN s_7_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_7(252) WHEN s_7_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_7(253) WHEN s_7_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_7(254) WHEN s_7_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_7(255);

  
  out0_160 <= gmul3_7(0) WHEN s_4_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_7(1) WHEN s_4_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_7(2) WHEN s_4_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_7(3) WHEN s_4_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_7(4) WHEN s_4_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_7(5) WHEN s_4_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_7(6) WHEN s_4_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_7(7) WHEN s_4_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_7(8) WHEN s_4_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_7(9) WHEN s_4_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_7(10) WHEN s_4_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_7(11) WHEN s_4_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_7(12) WHEN s_4_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_7(13) WHEN s_4_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_7(14) WHEN s_4_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_7(15) WHEN s_4_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_7(16) WHEN s_4_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_7(17) WHEN s_4_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_7(18) WHEN s_4_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_7(19) WHEN s_4_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_7(20) WHEN s_4_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_7(21) WHEN s_4_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_7(22) WHEN s_4_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_7(23) WHEN s_4_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_7(24) WHEN s_4_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_7(25) WHEN s_4_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_7(26) WHEN s_4_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_7(27) WHEN s_4_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_7(28) WHEN s_4_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_7(29) WHEN s_4_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_7(30) WHEN s_4_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_7(31) WHEN s_4_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_7(32) WHEN s_4_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_7(33) WHEN s_4_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_7(34) WHEN s_4_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_7(35) WHEN s_4_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_7(36) WHEN s_4_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_7(37) WHEN s_4_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_7(38) WHEN s_4_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_7(39) WHEN s_4_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_7(40) WHEN s_4_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_7(41) WHEN s_4_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_7(42) WHEN s_4_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_7(43) WHEN s_4_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_7(44) WHEN s_4_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_7(45) WHEN s_4_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_7(46) WHEN s_4_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_7(47) WHEN s_4_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_7(48) WHEN s_4_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_7(49) WHEN s_4_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_7(50) WHEN s_4_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_7(51) WHEN s_4_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_7(52) WHEN s_4_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_7(53) WHEN s_4_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_7(54) WHEN s_4_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_7(55) WHEN s_4_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_7(56) WHEN s_4_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_7(57) WHEN s_4_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_7(58) WHEN s_4_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_7(59) WHEN s_4_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_7(60) WHEN s_4_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_7(61) WHEN s_4_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_7(62) WHEN s_4_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_7(63) WHEN s_4_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_7(64) WHEN s_4_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_7(65) WHEN s_4_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_7(66) WHEN s_4_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_7(67) WHEN s_4_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_7(68) WHEN s_4_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_7(69) WHEN s_4_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_7(70) WHEN s_4_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_7(71) WHEN s_4_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_7(72) WHEN s_4_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_7(73) WHEN s_4_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_7(74) WHEN s_4_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_7(75) WHEN s_4_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_7(76) WHEN s_4_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_7(77) WHEN s_4_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_7(78) WHEN s_4_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_7(79) WHEN s_4_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_7(80) WHEN s_4_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_7(81) WHEN s_4_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_7(82) WHEN s_4_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_7(83) WHEN s_4_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_7(84) WHEN s_4_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_7(85) WHEN s_4_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_7(86) WHEN s_4_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_7(87) WHEN s_4_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_7(88) WHEN s_4_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_7(89) WHEN s_4_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_7(90) WHEN s_4_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_7(91) WHEN s_4_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_7(92) WHEN s_4_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_7(93) WHEN s_4_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_7(94) WHEN s_4_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_7(95) WHEN s_4_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_7(96) WHEN s_4_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_7(97) WHEN s_4_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_7(98) WHEN s_4_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_7(99) WHEN s_4_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_7(100) WHEN s_4_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_7(101) WHEN s_4_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_7(102) WHEN s_4_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_7(103) WHEN s_4_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_7(104) WHEN s_4_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_7(105) WHEN s_4_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_7(106) WHEN s_4_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_7(107) WHEN s_4_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_7(108) WHEN s_4_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_7(109) WHEN s_4_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_7(110) WHEN s_4_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_7(111) WHEN s_4_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_7(112) WHEN s_4_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_7(113) WHEN s_4_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_7(114) WHEN s_4_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_7(115) WHEN s_4_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_7(116) WHEN s_4_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_7(117) WHEN s_4_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_7(118) WHEN s_4_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_7(119) WHEN s_4_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_7(120) WHEN s_4_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_7(121) WHEN s_4_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_7(122) WHEN s_4_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_7(123) WHEN s_4_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_7(124) WHEN s_4_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_7(125) WHEN s_4_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_7(126) WHEN s_4_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_7(127) WHEN s_4_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_7(128) WHEN s_4_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_7(129) WHEN s_4_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_7(130) WHEN s_4_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_7(131) WHEN s_4_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_7(132) WHEN s_4_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_7(133) WHEN s_4_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_7(134) WHEN s_4_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_7(135) WHEN s_4_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_7(136) WHEN s_4_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_7(137) WHEN s_4_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_7(138) WHEN s_4_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_7(139) WHEN s_4_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_7(140) WHEN s_4_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_7(141) WHEN s_4_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_7(142) WHEN s_4_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_7(143) WHEN s_4_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_7(144) WHEN s_4_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_7(145) WHEN s_4_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_7(146) WHEN s_4_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_7(147) WHEN s_4_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_7(148) WHEN s_4_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_7(149) WHEN s_4_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_7(150) WHEN s_4_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_7(151) WHEN s_4_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_7(152) WHEN s_4_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_7(153) WHEN s_4_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_7(154) WHEN s_4_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_7(155) WHEN s_4_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_7(156) WHEN s_4_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_7(157) WHEN s_4_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_7(158) WHEN s_4_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_7(159) WHEN s_4_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_7(160) WHEN s_4_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_7(161) WHEN s_4_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_7(162) WHEN s_4_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_7(163) WHEN s_4_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_7(164) WHEN s_4_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_7(165) WHEN s_4_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_7(166) WHEN s_4_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_7(167) WHEN s_4_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_7(168) WHEN s_4_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_7(169) WHEN s_4_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_7(170) WHEN s_4_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_7(171) WHEN s_4_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_7(172) WHEN s_4_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_7(173) WHEN s_4_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_7(174) WHEN s_4_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_7(175) WHEN s_4_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_7(176) WHEN s_4_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_7(177) WHEN s_4_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_7(178) WHEN s_4_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_7(179) WHEN s_4_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_7(180) WHEN s_4_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_7(181) WHEN s_4_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_7(182) WHEN s_4_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_7(183) WHEN s_4_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_7(184) WHEN s_4_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_7(185) WHEN s_4_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_7(186) WHEN s_4_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_7(187) WHEN s_4_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_7(188) WHEN s_4_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_7(189) WHEN s_4_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_7(190) WHEN s_4_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_7(191) WHEN s_4_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_7(192) WHEN s_4_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_7(193) WHEN s_4_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_7(194) WHEN s_4_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_7(195) WHEN s_4_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_7(196) WHEN s_4_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_7(197) WHEN s_4_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_7(198) WHEN s_4_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_7(199) WHEN s_4_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_7(200) WHEN s_4_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_7(201) WHEN s_4_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_7(202) WHEN s_4_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_7(203) WHEN s_4_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_7(204) WHEN s_4_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_7(205) WHEN s_4_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_7(206) WHEN s_4_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_7(207) WHEN s_4_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_7(208) WHEN s_4_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_7(209) WHEN s_4_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_7(210) WHEN s_4_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_7(211) WHEN s_4_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_7(212) WHEN s_4_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_7(213) WHEN s_4_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_7(214) WHEN s_4_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_7(215) WHEN s_4_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_7(216) WHEN s_4_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_7(217) WHEN s_4_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_7(218) WHEN s_4_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_7(219) WHEN s_4_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_7(220) WHEN s_4_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_7(221) WHEN s_4_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_7(222) WHEN s_4_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_7(223) WHEN s_4_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_7(224) WHEN s_4_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_7(225) WHEN s_4_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_7(226) WHEN s_4_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_7(227) WHEN s_4_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_7(228) WHEN s_4_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_7(229) WHEN s_4_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_7(230) WHEN s_4_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_7(231) WHEN s_4_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_7(232) WHEN s_4_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_7(233) WHEN s_4_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_7(234) WHEN s_4_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_7(235) WHEN s_4_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_7(236) WHEN s_4_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_7(237) WHEN s_4_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_7(238) WHEN s_4_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_7(239) WHEN s_4_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_7(240) WHEN s_4_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_7(241) WHEN s_4_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_7(242) WHEN s_4_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_7(243) WHEN s_4_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_7(244) WHEN s_4_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_7(245) WHEN s_4_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_7(246) WHEN s_4_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_7(247) WHEN s_4_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_7(248) WHEN s_4_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_7(249) WHEN s_4_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_7(250) WHEN s_4_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_7(251) WHEN s_4_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_7(252) WHEN s_4_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_7(253) WHEN s_4_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_7(254) WHEN s_4_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_7(255);

  out0_161 <= out0_160 XOR s_5_1;

  b4_2 <= out0_161 XOR s_6_1;

  out0_162 <= b4_2 XOR out0_159;

  
  out0_163 <= gmul3_6(0) WHEN s_7_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_6(1) WHEN s_7_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_6(2) WHEN s_7_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_6(3) WHEN s_7_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_6(4) WHEN s_7_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_6(5) WHEN s_7_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_6(6) WHEN s_7_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_6(7) WHEN s_7_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_6(8) WHEN s_7_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_6(9) WHEN s_7_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_6(10) WHEN s_7_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_6(11) WHEN s_7_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_6(12) WHEN s_7_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_6(13) WHEN s_7_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_6(14) WHEN s_7_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_6(15) WHEN s_7_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_6(16) WHEN s_7_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_6(17) WHEN s_7_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_6(18) WHEN s_7_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_6(19) WHEN s_7_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_6(20) WHEN s_7_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_6(21) WHEN s_7_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_6(22) WHEN s_7_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_6(23) WHEN s_7_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_6(24) WHEN s_7_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_6(25) WHEN s_7_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_6(26) WHEN s_7_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_6(27) WHEN s_7_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_6(28) WHEN s_7_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_6(29) WHEN s_7_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_6(30) WHEN s_7_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_6(31) WHEN s_7_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_6(32) WHEN s_7_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_6(33) WHEN s_7_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_6(34) WHEN s_7_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_6(35) WHEN s_7_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_6(36) WHEN s_7_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_6(37) WHEN s_7_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_6(38) WHEN s_7_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_6(39) WHEN s_7_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_6(40) WHEN s_7_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_6(41) WHEN s_7_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_6(42) WHEN s_7_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_6(43) WHEN s_7_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_6(44) WHEN s_7_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_6(45) WHEN s_7_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_6(46) WHEN s_7_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_6(47) WHEN s_7_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_6(48) WHEN s_7_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_6(49) WHEN s_7_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_6(50) WHEN s_7_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_6(51) WHEN s_7_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_6(52) WHEN s_7_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_6(53) WHEN s_7_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_6(54) WHEN s_7_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_6(55) WHEN s_7_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_6(56) WHEN s_7_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_6(57) WHEN s_7_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_6(58) WHEN s_7_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_6(59) WHEN s_7_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_6(60) WHEN s_7_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_6(61) WHEN s_7_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_6(62) WHEN s_7_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_6(63) WHEN s_7_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_6(64) WHEN s_7_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_6(65) WHEN s_7_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_6(66) WHEN s_7_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_6(67) WHEN s_7_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_6(68) WHEN s_7_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_6(69) WHEN s_7_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_6(70) WHEN s_7_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_6(71) WHEN s_7_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_6(72) WHEN s_7_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_6(73) WHEN s_7_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_6(74) WHEN s_7_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_6(75) WHEN s_7_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_6(76) WHEN s_7_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_6(77) WHEN s_7_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_6(78) WHEN s_7_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_6(79) WHEN s_7_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_6(80) WHEN s_7_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_6(81) WHEN s_7_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_6(82) WHEN s_7_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_6(83) WHEN s_7_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_6(84) WHEN s_7_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_6(85) WHEN s_7_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_6(86) WHEN s_7_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_6(87) WHEN s_7_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_6(88) WHEN s_7_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_6(89) WHEN s_7_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_6(90) WHEN s_7_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_6(91) WHEN s_7_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_6(92) WHEN s_7_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_6(93) WHEN s_7_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_6(94) WHEN s_7_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_6(95) WHEN s_7_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_6(96) WHEN s_7_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_6(97) WHEN s_7_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_6(98) WHEN s_7_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_6(99) WHEN s_7_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_6(100) WHEN s_7_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_6(101) WHEN s_7_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_6(102) WHEN s_7_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_6(103) WHEN s_7_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_6(104) WHEN s_7_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_6(105) WHEN s_7_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_6(106) WHEN s_7_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_6(107) WHEN s_7_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_6(108) WHEN s_7_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_6(109) WHEN s_7_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_6(110) WHEN s_7_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_6(111) WHEN s_7_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_6(112) WHEN s_7_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_6(113) WHEN s_7_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_6(114) WHEN s_7_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_6(115) WHEN s_7_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_6(116) WHEN s_7_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_6(117) WHEN s_7_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_6(118) WHEN s_7_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_6(119) WHEN s_7_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_6(120) WHEN s_7_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_6(121) WHEN s_7_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_6(122) WHEN s_7_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_6(123) WHEN s_7_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_6(124) WHEN s_7_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_6(125) WHEN s_7_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_6(126) WHEN s_7_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_6(127) WHEN s_7_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_6(128) WHEN s_7_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_6(129) WHEN s_7_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_6(130) WHEN s_7_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_6(131) WHEN s_7_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_6(132) WHEN s_7_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_6(133) WHEN s_7_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_6(134) WHEN s_7_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_6(135) WHEN s_7_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_6(136) WHEN s_7_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_6(137) WHEN s_7_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_6(138) WHEN s_7_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_6(139) WHEN s_7_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_6(140) WHEN s_7_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_6(141) WHEN s_7_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_6(142) WHEN s_7_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_6(143) WHEN s_7_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_6(144) WHEN s_7_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_6(145) WHEN s_7_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_6(146) WHEN s_7_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_6(147) WHEN s_7_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_6(148) WHEN s_7_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_6(149) WHEN s_7_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_6(150) WHEN s_7_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_6(151) WHEN s_7_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_6(152) WHEN s_7_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_6(153) WHEN s_7_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_6(154) WHEN s_7_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_6(155) WHEN s_7_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_6(156) WHEN s_7_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_6(157) WHEN s_7_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_6(158) WHEN s_7_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_6(159) WHEN s_7_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_6(160) WHEN s_7_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_6(161) WHEN s_7_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_6(162) WHEN s_7_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_6(163) WHEN s_7_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_6(164) WHEN s_7_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_6(165) WHEN s_7_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_6(166) WHEN s_7_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_6(167) WHEN s_7_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_6(168) WHEN s_7_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_6(169) WHEN s_7_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_6(170) WHEN s_7_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_6(171) WHEN s_7_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_6(172) WHEN s_7_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_6(173) WHEN s_7_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_6(174) WHEN s_7_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_6(175) WHEN s_7_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_6(176) WHEN s_7_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_6(177) WHEN s_7_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_6(178) WHEN s_7_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_6(179) WHEN s_7_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_6(180) WHEN s_7_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_6(181) WHEN s_7_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_6(182) WHEN s_7_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_6(183) WHEN s_7_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_6(184) WHEN s_7_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_6(185) WHEN s_7_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_6(186) WHEN s_7_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_6(187) WHEN s_7_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_6(188) WHEN s_7_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_6(189) WHEN s_7_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_6(190) WHEN s_7_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_6(191) WHEN s_7_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_6(192) WHEN s_7_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_6(193) WHEN s_7_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_6(194) WHEN s_7_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_6(195) WHEN s_7_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_6(196) WHEN s_7_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_6(197) WHEN s_7_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_6(198) WHEN s_7_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_6(199) WHEN s_7_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_6(200) WHEN s_7_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_6(201) WHEN s_7_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_6(202) WHEN s_7_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_6(203) WHEN s_7_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_6(204) WHEN s_7_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_6(205) WHEN s_7_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_6(206) WHEN s_7_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_6(207) WHEN s_7_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_6(208) WHEN s_7_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_6(209) WHEN s_7_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_6(210) WHEN s_7_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_6(211) WHEN s_7_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_6(212) WHEN s_7_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_6(213) WHEN s_7_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_6(214) WHEN s_7_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_6(215) WHEN s_7_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_6(216) WHEN s_7_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_6(217) WHEN s_7_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_6(218) WHEN s_7_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_6(219) WHEN s_7_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_6(220) WHEN s_7_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_6(221) WHEN s_7_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_6(222) WHEN s_7_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_6(223) WHEN s_7_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_6(224) WHEN s_7_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_6(225) WHEN s_7_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_6(226) WHEN s_7_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_6(227) WHEN s_7_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_6(228) WHEN s_7_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_6(229) WHEN s_7_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_6(230) WHEN s_7_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_6(231) WHEN s_7_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_6(232) WHEN s_7_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_6(233) WHEN s_7_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_6(234) WHEN s_7_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_6(235) WHEN s_7_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_6(236) WHEN s_7_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_6(237) WHEN s_7_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_6(238) WHEN s_7_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_6(239) WHEN s_7_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_6(240) WHEN s_7_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_6(241) WHEN s_7_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_6(242) WHEN s_7_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_6(243) WHEN s_7_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_6(244) WHEN s_7_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_6(245) WHEN s_7_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_6(246) WHEN s_7_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_6(247) WHEN s_7_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_6(248) WHEN s_7_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_6(249) WHEN s_7_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_6(250) WHEN s_7_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_6(251) WHEN s_7_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_6(252) WHEN s_7_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_6(253) WHEN s_7_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_6(254) WHEN s_7_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_6(255);

  
  out0_164 <= gmul2_6(0) WHEN s_6_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_6(1) WHEN s_6_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_6(2) WHEN s_6_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_6(3) WHEN s_6_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_6(4) WHEN s_6_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_6(5) WHEN s_6_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_6(6) WHEN s_6_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_6(7) WHEN s_6_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_6(8) WHEN s_6_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_6(9) WHEN s_6_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_6(10) WHEN s_6_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_6(11) WHEN s_6_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_6(12) WHEN s_6_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_6(13) WHEN s_6_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_6(14) WHEN s_6_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_6(15) WHEN s_6_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_6(16) WHEN s_6_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_6(17) WHEN s_6_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_6(18) WHEN s_6_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_6(19) WHEN s_6_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_6(20) WHEN s_6_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_6(21) WHEN s_6_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_6(22) WHEN s_6_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_6(23) WHEN s_6_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_6(24) WHEN s_6_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_6(25) WHEN s_6_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_6(26) WHEN s_6_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_6(27) WHEN s_6_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_6(28) WHEN s_6_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_6(29) WHEN s_6_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_6(30) WHEN s_6_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_6(31) WHEN s_6_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_6(32) WHEN s_6_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_6(33) WHEN s_6_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_6(34) WHEN s_6_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_6(35) WHEN s_6_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_6(36) WHEN s_6_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_6(37) WHEN s_6_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_6(38) WHEN s_6_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_6(39) WHEN s_6_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_6(40) WHEN s_6_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_6(41) WHEN s_6_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_6(42) WHEN s_6_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_6(43) WHEN s_6_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_6(44) WHEN s_6_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_6(45) WHEN s_6_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_6(46) WHEN s_6_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_6(47) WHEN s_6_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_6(48) WHEN s_6_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_6(49) WHEN s_6_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_6(50) WHEN s_6_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_6(51) WHEN s_6_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_6(52) WHEN s_6_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_6(53) WHEN s_6_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_6(54) WHEN s_6_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_6(55) WHEN s_6_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_6(56) WHEN s_6_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_6(57) WHEN s_6_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_6(58) WHEN s_6_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_6(59) WHEN s_6_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_6(60) WHEN s_6_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_6(61) WHEN s_6_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_6(62) WHEN s_6_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_6(63) WHEN s_6_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_6(64) WHEN s_6_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_6(65) WHEN s_6_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_6(66) WHEN s_6_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_6(67) WHEN s_6_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_6(68) WHEN s_6_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_6(69) WHEN s_6_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_6(70) WHEN s_6_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_6(71) WHEN s_6_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_6(72) WHEN s_6_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_6(73) WHEN s_6_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_6(74) WHEN s_6_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_6(75) WHEN s_6_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_6(76) WHEN s_6_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_6(77) WHEN s_6_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_6(78) WHEN s_6_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_6(79) WHEN s_6_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_6(80) WHEN s_6_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_6(81) WHEN s_6_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_6(82) WHEN s_6_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_6(83) WHEN s_6_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_6(84) WHEN s_6_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_6(85) WHEN s_6_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_6(86) WHEN s_6_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_6(87) WHEN s_6_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_6(88) WHEN s_6_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_6(89) WHEN s_6_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_6(90) WHEN s_6_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_6(91) WHEN s_6_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_6(92) WHEN s_6_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_6(93) WHEN s_6_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_6(94) WHEN s_6_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_6(95) WHEN s_6_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_6(96) WHEN s_6_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_6(97) WHEN s_6_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_6(98) WHEN s_6_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_6(99) WHEN s_6_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_6(100) WHEN s_6_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_6(101) WHEN s_6_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_6(102) WHEN s_6_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_6(103) WHEN s_6_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_6(104) WHEN s_6_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_6(105) WHEN s_6_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_6(106) WHEN s_6_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_6(107) WHEN s_6_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_6(108) WHEN s_6_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_6(109) WHEN s_6_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_6(110) WHEN s_6_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_6(111) WHEN s_6_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_6(112) WHEN s_6_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_6(113) WHEN s_6_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_6(114) WHEN s_6_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_6(115) WHEN s_6_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_6(116) WHEN s_6_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_6(117) WHEN s_6_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_6(118) WHEN s_6_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_6(119) WHEN s_6_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_6(120) WHEN s_6_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_6(121) WHEN s_6_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_6(122) WHEN s_6_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_6(123) WHEN s_6_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_6(124) WHEN s_6_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_6(125) WHEN s_6_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_6(126) WHEN s_6_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_6(127) WHEN s_6_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_6(128) WHEN s_6_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_6(129) WHEN s_6_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_6(130) WHEN s_6_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_6(131) WHEN s_6_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_6(132) WHEN s_6_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_6(133) WHEN s_6_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_6(134) WHEN s_6_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_6(135) WHEN s_6_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_6(136) WHEN s_6_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_6(137) WHEN s_6_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_6(138) WHEN s_6_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_6(139) WHEN s_6_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_6(140) WHEN s_6_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_6(141) WHEN s_6_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_6(142) WHEN s_6_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_6(143) WHEN s_6_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_6(144) WHEN s_6_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_6(145) WHEN s_6_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_6(146) WHEN s_6_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_6(147) WHEN s_6_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_6(148) WHEN s_6_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_6(149) WHEN s_6_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_6(150) WHEN s_6_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_6(151) WHEN s_6_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_6(152) WHEN s_6_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_6(153) WHEN s_6_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_6(154) WHEN s_6_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_6(155) WHEN s_6_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_6(156) WHEN s_6_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_6(157) WHEN s_6_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_6(158) WHEN s_6_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_6(159) WHEN s_6_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_6(160) WHEN s_6_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_6(161) WHEN s_6_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_6(162) WHEN s_6_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_6(163) WHEN s_6_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_6(164) WHEN s_6_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_6(165) WHEN s_6_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_6(166) WHEN s_6_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_6(167) WHEN s_6_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_6(168) WHEN s_6_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_6(169) WHEN s_6_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_6(170) WHEN s_6_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_6(171) WHEN s_6_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_6(172) WHEN s_6_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_6(173) WHEN s_6_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_6(174) WHEN s_6_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_6(175) WHEN s_6_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_6(176) WHEN s_6_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_6(177) WHEN s_6_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_6(178) WHEN s_6_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_6(179) WHEN s_6_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_6(180) WHEN s_6_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_6(181) WHEN s_6_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_6(182) WHEN s_6_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_6(183) WHEN s_6_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_6(184) WHEN s_6_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_6(185) WHEN s_6_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_6(186) WHEN s_6_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_6(187) WHEN s_6_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_6(188) WHEN s_6_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_6(189) WHEN s_6_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_6(190) WHEN s_6_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_6(191) WHEN s_6_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_6(192) WHEN s_6_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_6(193) WHEN s_6_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_6(194) WHEN s_6_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_6(195) WHEN s_6_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_6(196) WHEN s_6_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_6(197) WHEN s_6_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_6(198) WHEN s_6_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_6(199) WHEN s_6_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_6(200) WHEN s_6_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_6(201) WHEN s_6_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_6(202) WHEN s_6_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_6(203) WHEN s_6_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_6(204) WHEN s_6_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_6(205) WHEN s_6_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_6(206) WHEN s_6_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_6(207) WHEN s_6_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_6(208) WHEN s_6_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_6(209) WHEN s_6_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_6(210) WHEN s_6_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_6(211) WHEN s_6_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_6(212) WHEN s_6_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_6(213) WHEN s_6_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_6(214) WHEN s_6_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_6(215) WHEN s_6_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_6(216) WHEN s_6_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_6(217) WHEN s_6_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_6(218) WHEN s_6_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_6(219) WHEN s_6_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_6(220) WHEN s_6_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_6(221) WHEN s_6_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_6(222) WHEN s_6_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_6(223) WHEN s_6_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_6(224) WHEN s_6_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_6(225) WHEN s_6_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_6(226) WHEN s_6_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_6(227) WHEN s_6_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_6(228) WHEN s_6_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_6(229) WHEN s_6_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_6(230) WHEN s_6_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_6(231) WHEN s_6_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_6(232) WHEN s_6_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_6(233) WHEN s_6_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_6(234) WHEN s_6_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_6(235) WHEN s_6_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_6(236) WHEN s_6_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_6(237) WHEN s_6_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_6(238) WHEN s_6_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_6(239) WHEN s_6_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_6(240) WHEN s_6_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_6(241) WHEN s_6_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_6(242) WHEN s_6_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_6(243) WHEN s_6_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_6(244) WHEN s_6_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_6(245) WHEN s_6_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_6(246) WHEN s_6_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_6(247) WHEN s_6_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_6(248) WHEN s_6_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_6(249) WHEN s_6_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_6(250) WHEN s_6_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_6(251) WHEN s_6_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_6(252) WHEN s_6_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_6(253) WHEN s_6_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_6(254) WHEN s_6_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_6(255);

  out0_165 <= s_4_1 XOR s_5_1;

  b3_2 <= out0_165 XOR out0_164;

  out0_166 <= b3_2 XOR out0_163;

  
  out0_167 <= gmul3_5(0) WHEN s_6_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_5(1) WHEN s_6_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_5(2) WHEN s_6_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_5(3) WHEN s_6_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_5(4) WHEN s_6_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_5(5) WHEN s_6_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_5(6) WHEN s_6_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_5(7) WHEN s_6_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_5(8) WHEN s_6_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_5(9) WHEN s_6_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_5(10) WHEN s_6_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_5(11) WHEN s_6_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_5(12) WHEN s_6_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_5(13) WHEN s_6_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_5(14) WHEN s_6_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_5(15) WHEN s_6_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_5(16) WHEN s_6_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_5(17) WHEN s_6_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_5(18) WHEN s_6_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_5(19) WHEN s_6_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_5(20) WHEN s_6_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_5(21) WHEN s_6_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_5(22) WHEN s_6_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_5(23) WHEN s_6_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_5(24) WHEN s_6_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_5(25) WHEN s_6_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_5(26) WHEN s_6_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_5(27) WHEN s_6_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_5(28) WHEN s_6_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_5(29) WHEN s_6_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_5(30) WHEN s_6_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_5(31) WHEN s_6_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_5(32) WHEN s_6_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_5(33) WHEN s_6_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_5(34) WHEN s_6_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_5(35) WHEN s_6_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_5(36) WHEN s_6_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_5(37) WHEN s_6_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_5(38) WHEN s_6_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_5(39) WHEN s_6_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_5(40) WHEN s_6_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_5(41) WHEN s_6_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_5(42) WHEN s_6_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_5(43) WHEN s_6_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_5(44) WHEN s_6_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_5(45) WHEN s_6_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_5(46) WHEN s_6_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_5(47) WHEN s_6_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_5(48) WHEN s_6_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_5(49) WHEN s_6_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_5(50) WHEN s_6_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_5(51) WHEN s_6_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_5(52) WHEN s_6_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_5(53) WHEN s_6_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_5(54) WHEN s_6_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_5(55) WHEN s_6_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_5(56) WHEN s_6_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_5(57) WHEN s_6_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_5(58) WHEN s_6_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_5(59) WHEN s_6_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_5(60) WHEN s_6_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_5(61) WHEN s_6_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_5(62) WHEN s_6_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_5(63) WHEN s_6_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_5(64) WHEN s_6_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_5(65) WHEN s_6_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_5(66) WHEN s_6_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_5(67) WHEN s_6_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_5(68) WHEN s_6_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_5(69) WHEN s_6_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_5(70) WHEN s_6_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_5(71) WHEN s_6_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_5(72) WHEN s_6_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_5(73) WHEN s_6_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_5(74) WHEN s_6_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_5(75) WHEN s_6_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_5(76) WHEN s_6_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_5(77) WHEN s_6_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_5(78) WHEN s_6_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_5(79) WHEN s_6_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_5(80) WHEN s_6_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_5(81) WHEN s_6_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_5(82) WHEN s_6_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_5(83) WHEN s_6_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_5(84) WHEN s_6_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_5(85) WHEN s_6_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_5(86) WHEN s_6_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_5(87) WHEN s_6_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_5(88) WHEN s_6_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_5(89) WHEN s_6_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_5(90) WHEN s_6_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_5(91) WHEN s_6_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_5(92) WHEN s_6_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_5(93) WHEN s_6_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_5(94) WHEN s_6_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_5(95) WHEN s_6_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_5(96) WHEN s_6_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_5(97) WHEN s_6_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_5(98) WHEN s_6_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_5(99) WHEN s_6_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_5(100) WHEN s_6_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_5(101) WHEN s_6_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_5(102) WHEN s_6_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_5(103) WHEN s_6_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_5(104) WHEN s_6_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_5(105) WHEN s_6_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_5(106) WHEN s_6_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_5(107) WHEN s_6_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_5(108) WHEN s_6_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_5(109) WHEN s_6_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_5(110) WHEN s_6_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_5(111) WHEN s_6_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_5(112) WHEN s_6_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_5(113) WHEN s_6_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_5(114) WHEN s_6_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_5(115) WHEN s_6_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_5(116) WHEN s_6_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_5(117) WHEN s_6_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_5(118) WHEN s_6_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_5(119) WHEN s_6_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_5(120) WHEN s_6_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_5(121) WHEN s_6_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_5(122) WHEN s_6_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_5(123) WHEN s_6_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_5(124) WHEN s_6_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_5(125) WHEN s_6_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_5(126) WHEN s_6_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_5(127) WHEN s_6_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_5(128) WHEN s_6_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_5(129) WHEN s_6_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_5(130) WHEN s_6_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_5(131) WHEN s_6_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_5(132) WHEN s_6_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_5(133) WHEN s_6_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_5(134) WHEN s_6_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_5(135) WHEN s_6_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_5(136) WHEN s_6_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_5(137) WHEN s_6_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_5(138) WHEN s_6_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_5(139) WHEN s_6_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_5(140) WHEN s_6_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_5(141) WHEN s_6_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_5(142) WHEN s_6_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_5(143) WHEN s_6_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_5(144) WHEN s_6_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_5(145) WHEN s_6_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_5(146) WHEN s_6_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_5(147) WHEN s_6_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_5(148) WHEN s_6_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_5(149) WHEN s_6_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_5(150) WHEN s_6_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_5(151) WHEN s_6_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_5(152) WHEN s_6_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_5(153) WHEN s_6_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_5(154) WHEN s_6_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_5(155) WHEN s_6_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_5(156) WHEN s_6_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_5(157) WHEN s_6_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_5(158) WHEN s_6_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_5(159) WHEN s_6_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_5(160) WHEN s_6_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_5(161) WHEN s_6_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_5(162) WHEN s_6_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_5(163) WHEN s_6_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_5(164) WHEN s_6_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_5(165) WHEN s_6_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_5(166) WHEN s_6_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_5(167) WHEN s_6_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_5(168) WHEN s_6_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_5(169) WHEN s_6_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_5(170) WHEN s_6_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_5(171) WHEN s_6_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_5(172) WHEN s_6_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_5(173) WHEN s_6_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_5(174) WHEN s_6_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_5(175) WHEN s_6_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_5(176) WHEN s_6_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_5(177) WHEN s_6_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_5(178) WHEN s_6_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_5(179) WHEN s_6_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_5(180) WHEN s_6_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_5(181) WHEN s_6_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_5(182) WHEN s_6_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_5(183) WHEN s_6_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_5(184) WHEN s_6_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_5(185) WHEN s_6_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_5(186) WHEN s_6_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_5(187) WHEN s_6_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_5(188) WHEN s_6_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_5(189) WHEN s_6_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_5(190) WHEN s_6_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_5(191) WHEN s_6_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_5(192) WHEN s_6_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_5(193) WHEN s_6_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_5(194) WHEN s_6_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_5(195) WHEN s_6_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_5(196) WHEN s_6_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_5(197) WHEN s_6_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_5(198) WHEN s_6_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_5(199) WHEN s_6_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_5(200) WHEN s_6_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_5(201) WHEN s_6_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_5(202) WHEN s_6_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_5(203) WHEN s_6_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_5(204) WHEN s_6_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_5(205) WHEN s_6_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_5(206) WHEN s_6_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_5(207) WHEN s_6_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_5(208) WHEN s_6_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_5(209) WHEN s_6_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_5(210) WHEN s_6_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_5(211) WHEN s_6_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_5(212) WHEN s_6_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_5(213) WHEN s_6_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_5(214) WHEN s_6_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_5(215) WHEN s_6_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_5(216) WHEN s_6_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_5(217) WHEN s_6_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_5(218) WHEN s_6_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_5(219) WHEN s_6_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_5(220) WHEN s_6_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_5(221) WHEN s_6_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_5(222) WHEN s_6_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_5(223) WHEN s_6_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_5(224) WHEN s_6_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_5(225) WHEN s_6_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_5(226) WHEN s_6_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_5(227) WHEN s_6_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_5(228) WHEN s_6_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_5(229) WHEN s_6_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_5(230) WHEN s_6_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_5(231) WHEN s_6_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_5(232) WHEN s_6_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_5(233) WHEN s_6_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_5(234) WHEN s_6_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_5(235) WHEN s_6_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_5(236) WHEN s_6_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_5(237) WHEN s_6_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_5(238) WHEN s_6_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_5(239) WHEN s_6_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_5(240) WHEN s_6_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_5(241) WHEN s_6_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_5(242) WHEN s_6_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_5(243) WHEN s_6_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_5(244) WHEN s_6_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_5(245) WHEN s_6_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_5(246) WHEN s_6_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_5(247) WHEN s_6_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_5(248) WHEN s_6_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_5(249) WHEN s_6_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_5(250) WHEN s_6_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_5(251) WHEN s_6_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_5(252) WHEN s_6_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_5(253) WHEN s_6_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_5(254) WHEN s_6_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_5(255);

  
  out0_168 <= gmul2_5(0) WHEN s_5_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_5(1) WHEN s_5_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_5(2) WHEN s_5_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_5(3) WHEN s_5_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_5(4) WHEN s_5_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_5(5) WHEN s_5_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_5(6) WHEN s_5_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_5(7) WHEN s_5_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_5(8) WHEN s_5_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_5(9) WHEN s_5_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_5(10) WHEN s_5_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_5(11) WHEN s_5_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_5(12) WHEN s_5_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_5(13) WHEN s_5_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_5(14) WHEN s_5_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_5(15) WHEN s_5_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_5(16) WHEN s_5_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_5(17) WHEN s_5_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_5(18) WHEN s_5_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_5(19) WHEN s_5_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_5(20) WHEN s_5_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_5(21) WHEN s_5_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_5(22) WHEN s_5_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_5(23) WHEN s_5_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_5(24) WHEN s_5_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_5(25) WHEN s_5_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_5(26) WHEN s_5_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_5(27) WHEN s_5_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_5(28) WHEN s_5_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_5(29) WHEN s_5_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_5(30) WHEN s_5_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_5(31) WHEN s_5_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_5(32) WHEN s_5_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_5(33) WHEN s_5_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_5(34) WHEN s_5_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_5(35) WHEN s_5_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_5(36) WHEN s_5_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_5(37) WHEN s_5_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_5(38) WHEN s_5_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_5(39) WHEN s_5_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_5(40) WHEN s_5_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_5(41) WHEN s_5_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_5(42) WHEN s_5_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_5(43) WHEN s_5_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_5(44) WHEN s_5_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_5(45) WHEN s_5_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_5(46) WHEN s_5_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_5(47) WHEN s_5_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_5(48) WHEN s_5_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_5(49) WHEN s_5_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_5(50) WHEN s_5_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_5(51) WHEN s_5_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_5(52) WHEN s_5_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_5(53) WHEN s_5_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_5(54) WHEN s_5_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_5(55) WHEN s_5_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_5(56) WHEN s_5_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_5(57) WHEN s_5_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_5(58) WHEN s_5_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_5(59) WHEN s_5_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_5(60) WHEN s_5_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_5(61) WHEN s_5_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_5(62) WHEN s_5_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_5(63) WHEN s_5_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_5(64) WHEN s_5_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_5(65) WHEN s_5_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_5(66) WHEN s_5_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_5(67) WHEN s_5_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_5(68) WHEN s_5_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_5(69) WHEN s_5_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_5(70) WHEN s_5_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_5(71) WHEN s_5_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_5(72) WHEN s_5_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_5(73) WHEN s_5_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_5(74) WHEN s_5_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_5(75) WHEN s_5_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_5(76) WHEN s_5_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_5(77) WHEN s_5_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_5(78) WHEN s_5_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_5(79) WHEN s_5_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_5(80) WHEN s_5_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_5(81) WHEN s_5_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_5(82) WHEN s_5_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_5(83) WHEN s_5_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_5(84) WHEN s_5_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_5(85) WHEN s_5_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_5(86) WHEN s_5_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_5(87) WHEN s_5_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_5(88) WHEN s_5_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_5(89) WHEN s_5_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_5(90) WHEN s_5_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_5(91) WHEN s_5_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_5(92) WHEN s_5_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_5(93) WHEN s_5_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_5(94) WHEN s_5_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_5(95) WHEN s_5_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_5(96) WHEN s_5_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_5(97) WHEN s_5_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_5(98) WHEN s_5_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_5(99) WHEN s_5_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_5(100) WHEN s_5_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_5(101) WHEN s_5_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_5(102) WHEN s_5_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_5(103) WHEN s_5_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_5(104) WHEN s_5_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_5(105) WHEN s_5_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_5(106) WHEN s_5_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_5(107) WHEN s_5_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_5(108) WHEN s_5_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_5(109) WHEN s_5_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_5(110) WHEN s_5_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_5(111) WHEN s_5_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_5(112) WHEN s_5_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_5(113) WHEN s_5_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_5(114) WHEN s_5_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_5(115) WHEN s_5_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_5(116) WHEN s_5_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_5(117) WHEN s_5_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_5(118) WHEN s_5_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_5(119) WHEN s_5_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_5(120) WHEN s_5_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_5(121) WHEN s_5_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_5(122) WHEN s_5_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_5(123) WHEN s_5_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_5(124) WHEN s_5_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_5(125) WHEN s_5_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_5(126) WHEN s_5_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_5(127) WHEN s_5_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_5(128) WHEN s_5_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_5(129) WHEN s_5_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_5(130) WHEN s_5_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_5(131) WHEN s_5_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_5(132) WHEN s_5_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_5(133) WHEN s_5_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_5(134) WHEN s_5_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_5(135) WHEN s_5_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_5(136) WHEN s_5_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_5(137) WHEN s_5_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_5(138) WHEN s_5_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_5(139) WHEN s_5_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_5(140) WHEN s_5_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_5(141) WHEN s_5_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_5(142) WHEN s_5_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_5(143) WHEN s_5_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_5(144) WHEN s_5_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_5(145) WHEN s_5_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_5(146) WHEN s_5_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_5(147) WHEN s_5_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_5(148) WHEN s_5_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_5(149) WHEN s_5_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_5(150) WHEN s_5_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_5(151) WHEN s_5_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_5(152) WHEN s_5_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_5(153) WHEN s_5_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_5(154) WHEN s_5_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_5(155) WHEN s_5_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_5(156) WHEN s_5_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_5(157) WHEN s_5_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_5(158) WHEN s_5_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_5(159) WHEN s_5_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_5(160) WHEN s_5_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_5(161) WHEN s_5_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_5(162) WHEN s_5_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_5(163) WHEN s_5_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_5(164) WHEN s_5_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_5(165) WHEN s_5_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_5(166) WHEN s_5_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_5(167) WHEN s_5_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_5(168) WHEN s_5_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_5(169) WHEN s_5_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_5(170) WHEN s_5_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_5(171) WHEN s_5_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_5(172) WHEN s_5_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_5(173) WHEN s_5_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_5(174) WHEN s_5_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_5(175) WHEN s_5_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_5(176) WHEN s_5_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_5(177) WHEN s_5_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_5(178) WHEN s_5_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_5(179) WHEN s_5_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_5(180) WHEN s_5_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_5(181) WHEN s_5_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_5(182) WHEN s_5_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_5(183) WHEN s_5_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_5(184) WHEN s_5_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_5(185) WHEN s_5_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_5(186) WHEN s_5_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_5(187) WHEN s_5_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_5(188) WHEN s_5_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_5(189) WHEN s_5_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_5(190) WHEN s_5_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_5(191) WHEN s_5_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_5(192) WHEN s_5_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_5(193) WHEN s_5_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_5(194) WHEN s_5_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_5(195) WHEN s_5_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_5(196) WHEN s_5_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_5(197) WHEN s_5_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_5(198) WHEN s_5_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_5(199) WHEN s_5_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_5(200) WHEN s_5_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_5(201) WHEN s_5_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_5(202) WHEN s_5_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_5(203) WHEN s_5_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_5(204) WHEN s_5_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_5(205) WHEN s_5_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_5(206) WHEN s_5_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_5(207) WHEN s_5_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_5(208) WHEN s_5_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_5(209) WHEN s_5_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_5(210) WHEN s_5_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_5(211) WHEN s_5_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_5(212) WHEN s_5_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_5(213) WHEN s_5_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_5(214) WHEN s_5_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_5(215) WHEN s_5_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_5(216) WHEN s_5_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_5(217) WHEN s_5_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_5(218) WHEN s_5_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_5(219) WHEN s_5_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_5(220) WHEN s_5_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_5(221) WHEN s_5_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_5(222) WHEN s_5_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_5(223) WHEN s_5_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_5(224) WHEN s_5_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_5(225) WHEN s_5_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_5(226) WHEN s_5_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_5(227) WHEN s_5_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_5(228) WHEN s_5_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_5(229) WHEN s_5_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_5(230) WHEN s_5_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_5(231) WHEN s_5_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_5(232) WHEN s_5_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_5(233) WHEN s_5_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_5(234) WHEN s_5_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_5(235) WHEN s_5_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_5(236) WHEN s_5_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_5(237) WHEN s_5_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_5(238) WHEN s_5_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_5(239) WHEN s_5_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_5(240) WHEN s_5_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_5(241) WHEN s_5_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_5(242) WHEN s_5_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_5(243) WHEN s_5_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_5(244) WHEN s_5_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_5(245) WHEN s_5_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_5(246) WHEN s_5_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_5(247) WHEN s_5_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_5(248) WHEN s_5_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_5(249) WHEN s_5_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_5(250) WHEN s_5_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_5(251) WHEN s_5_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_5(252) WHEN s_5_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_5(253) WHEN s_5_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_5(254) WHEN s_5_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_5(255);

  out0_169 <= s_4_1 XOR out0_168;

  b2_2 <= out0_169 XOR out0_167;

  out0_170 <= b2_2 XOR s_7_1;

  s_7_1 <= s_s_6(7);

  s_6_1 <= s_s_6(6);

  s_5_1 <= s_s_6(5);

  
  out0_171 <= gmul3_4(0) WHEN s_5_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_4(1) WHEN s_5_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_4(2) WHEN s_5_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_4(3) WHEN s_5_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_4(4) WHEN s_5_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_4(5) WHEN s_5_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_4(6) WHEN s_5_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_4(7) WHEN s_5_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_4(8) WHEN s_5_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_4(9) WHEN s_5_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_4(10) WHEN s_5_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_4(11) WHEN s_5_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_4(12) WHEN s_5_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_4(13) WHEN s_5_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_4(14) WHEN s_5_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_4(15) WHEN s_5_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_4(16) WHEN s_5_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_4(17) WHEN s_5_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_4(18) WHEN s_5_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_4(19) WHEN s_5_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_4(20) WHEN s_5_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_4(21) WHEN s_5_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_4(22) WHEN s_5_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_4(23) WHEN s_5_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_4(24) WHEN s_5_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_4(25) WHEN s_5_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_4(26) WHEN s_5_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_4(27) WHEN s_5_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_4(28) WHEN s_5_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_4(29) WHEN s_5_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_4(30) WHEN s_5_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_4(31) WHEN s_5_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_4(32) WHEN s_5_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_4(33) WHEN s_5_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_4(34) WHEN s_5_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_4(35) WHEN s_5_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_4(36) WHEN s_5_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_4(37) WHEN s_5_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_4(38) WHEN s_5_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_4(39) WHEN s_5_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_4(40) WHEN s_5_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_4(41) WHEN s_5_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_4(42) WHEN s_5_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_4(43) WHEN s_5_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_4(44) WHEN s_5_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_4(45) WHEN s_5_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_4(46) WHEN s_5_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_4(47) WHEN s_5_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_4(48) WHEN s_5_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_4(49) WHEN s_5_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_4(50) WHEN s_5_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_4(51) WHEN s_5_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_4(52) WHEN s_5_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_4(53) WHEN s_5_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_4(54) WHEN s_5_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_4(55) WHEN s_5_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_4(56) WHEN s_5_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_4(57) WHEN s_5_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_4(58) WHEN s_5_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_4(59) WHEN s_5_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_4(60) WHEN s_5_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_4(61) WHEN s_5_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_4(62) WHEN s_5_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_4(63) WHEN s_5_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_4(64) WHEN s_5_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_4(65) WHEN s_5_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_4(66) WHEN s_5_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_4(67) WHEN s_5_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_4(68) WHEN s_5_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_4(69) WHEN s_5_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_4(70) WHEN s_5_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_4(71) WHEN s_5_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_4(72) WHEN s_5_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_4(73) WHEN s_5_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_4(74) WHEN s_5_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_4(75) WHEN s_5_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_4(76) WHEN s_5_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_4(77) WHEN s_5_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_4(78) WHEN s_5_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_4(79) WHEN s_5_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_4(80) WHEN s_5_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_4(81) WHEN s_5_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_4(82) WHEN s_5_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_4(83) WHEN s_5_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_4(84) WHEN s_5_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_4(85) WHEN s_5_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_4(86) WHEN s_5_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_4(87) WHEN s_5_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_4(88) WHEN s_5_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_4(89) WHEN s_5_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_4(90) WHEN s_5_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_4(91) WHEN s_5_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_4(92) WHEN s_5_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_4(93) WHEN s_5_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_4(94) WHEN s_5_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_4(95) WHEN s_5_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_4(96) WHEN s_5_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_4(97) WHEN s_5_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_4(98) WHEN s_5_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_4(99) WHEN s_5_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_4(100) WHEN s_5_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_4(101) WHEN s_5_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_4(102) WHEN s_5_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_4(103) WHEN s_5_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_4(104) WHEN s_5_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_4(105) WHEN s_5_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_4(106) WHEN s_5_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_4(107) WHEN s_5_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_4(108) WHEN s_5_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_4(109) WHEN s_5_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_4(110) WHEN s_5_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_4(111) WHEN s_5_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_4(112) WHEN s_5_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_4(113) WHEN s_5_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_4(114) WHEN s_5_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_4(115) WHEN s_5_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_4(116) WHEN s_5_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_4(117) WHEN s_5_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_4(118) WHEN s_5_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_4(119) WHEN s_5_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_4(120) WHEN s_5_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_4(121) WHEN s_5_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_4(122) WHEN s_5_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_4(123) WHEN s_5_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_4(124) WHEN s_5_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_4(125) WHEN s_5_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_4(126) WHEN s_5_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_4(127) WHEN s_5_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_4(128) WHEN s_5_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_4(129) WHEN s_5_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_4(130) WHEN s_5_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_4(131) WHEN s_5_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_4(132) WHEN s_5_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_4(133) WHEN s_5_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_4(134) WHEN s_5_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_4(135) WHEN s_5_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_4(136) WHEN s_5_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_4(137) WHEN s_5_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_4(138) WHEN s_5_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_4(139) WHEN s_5_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_4(140) WHEN s_5_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_4(141) WHEN s_5_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_4(142) WHEN s_5_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_4(143) WHEN s_5_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_4(144) WHEN s_5_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_4(145) WHEN s_5_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_4(146) WHEN s_5_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_4(147) WHEN s_5_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_4(148) WHEN s_5_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_4(149) WHEN s_5_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_4(150) WHEN s_5_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_4(151) WHEN s_5_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_4(152) WHEN s_5_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_4(153) WHEN s_5_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_4(154) WHEN s_5_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_4(155) WHEN s_5_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_4(156) WHEN s_5_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_4(157) WHEN s_5_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_4(158) WHEN s_5_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_4(159) WHEN s_5_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_4(160) WHEN s_5_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_4(161) WHEN s_5_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_4(162) WHEN s_5_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_4(163) WHEN s_5_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_4(164) WHEN s_5_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_4(165) WHEN s_5_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_4(166) WHEN s_5_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_4(167) WHEN s_5_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_4(168) WHEN s_5_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_4(169) WHEN s_5_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_4(170) WHEN s_5_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_4(171) WHEN s_5_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_4(172) WHEN s_5_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_4(173) WHEN s_5_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_4(174) WHEN s_5_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_4(175) WHEN s_5_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_4(176) WHEN s_5_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_4(177) WHEN s_5_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_4(178) WHEN s_5_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_4(179) WHEN s_5_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_4(180) WHEN s_5_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_4(181) WHEN s_5_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_4(182) WHEN s_5_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_4(183) WHEN s_5_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_4(184) WHEN s_5_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_4(185) WHEN s_5_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_4(186) WHEN s_5_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_4(187) WHEN s_5_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_4(188) WHEN s_5_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_4(189) WHEN s_5_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_4(190) WHEN s_5_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_4(191) WHEN s_5_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_4(192) WHEN s_5_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_4(193) WHEN s_5_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_4(194) WHEN s_5_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_4(195) WHEN s_5_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_4(196) WHEN s_5_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_4(197) WHEN s_5_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_4(198) WHEN s_5_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_4(199) WHEN s_5_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_4(200) WHEN s_5_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_4(201) WHEN s_5_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_4(202) WHEN s_5_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_4(203) WHEN s_5_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_4(204) WHEN s_5_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_4(205) WHEN s_5_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_4(206) WHEN s_5_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_4(207) WHEN s_5_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_4(208) WHEN s_5_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_4(209) WHEN s_5_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_4(210) WHEN s_5_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_4(211) WHEN s_5_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_4(212) WHEN s_5_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_4(213) WHEN s_5_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_4(214) WHEN s_5_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_4(215) WHEN s_5_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_4(216) WHEN s_5_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_4(217) WHEN s_5_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_4(218) WHEN s_5_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_4(219) WHEN s_5_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_4(220) WHEN s_5_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_4(221) WHEN s_5_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_4(222) WHEN s_5_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_4(223) WHEN s_5_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_4(224) WHEN s_5_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_4(225) WHEN s_5_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_4(226) WHEN s_5_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_4(227) WHEN s_5_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_4(228) WHEN s_5_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_4(229) WHEN s_5_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_4(230) WHEN s_5_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_4(231) WHEN s_5_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_4(232) WHEN s_5_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_4(233) WHEN s_5_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_4(234) WHEN s_5_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_4(235) WHEN s_5_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_4(236) WHEN s_5_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_4(237) WHEN s_5_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_4(238) WHEN s_5_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_4(239) WHEN s_5_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_4(240) WHEN s_5_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_4(241) WHEN s_5_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_4(242) WHEN s_5_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_4(243) WHEN s_5_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_4(244) WHEN s_5_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_4(245) WHEN s_5_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_4(246) WHEN s_5_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_4(247) WHEN s_5_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_4(248) WHEN s_5_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_4(249) WHEN s_5_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_4(250) WHEN s_5_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_4(251) WHEN s_5_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_4(252) WHEN s_5_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_4(253) WHEN s_5_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_4(254) WHEN s_5_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_4(255);

  s_4_1 <= s_s_6(4);

  
  out0_172 <= gmul2_4(0) WHEN s_4_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_4(1) WHEN s_4_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_4(2) WHEN s_4_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_4(3) WHEN s_4_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_4(4) WHEN s_4_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_4(5) WHEN s_4_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_4(6) WHEN s_4_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_4(7) WHEN s_4_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_4(8) WHEN s_4_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_4(9) WHEN s_4_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_4(10) WHEN s_4_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_4(11) WHEN s_4_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_4(12) WHEN s_4_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_4(13) WHEN s_4_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_4(14) WHEN s_4_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_4(15) WHEN s_4_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_4(16) WHEN s_4_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_4(17) WHEN s_4_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_4(18) WHEN s_4_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_4(19) WHEN s_4_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_4(20) WHEN s_4_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_4(21) WHEN s_4_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_4(22) WHEN s_4_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_4(23) WHEN s_4_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_4(24) WHEN s_4_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_4(25) WHEN s_4_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_4(26) WHEN s_4_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_4(27) WHEN s_4_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_4(28) WHEN s_4_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_4(29) WHEN s_4_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_4(30) WHEN s_4_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_4(31) WHEN s_4_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_4(32) WHEN s_4_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_4(33) WHEN s_4_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_4(34) WHEN s_4_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_4(35) WHEN s_4_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_4(36) WHEN s_4_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_4(37) WHEN s_4_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_4(38) WHEN s_4_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_4(39) WHEN s_4_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_4(40) WHEN s_4_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_4(41) WHEN s_4_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_4(42) WHEN s_4_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_4(43) WHEN s_4_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_4(44) WHEN s_4_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_4(45) WHEN s_4_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_4(46) WHEN s_4_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_4(47) WHEN s_4_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_4(48) WHEN s_4_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_4(49) WHEN s_4_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_4(50) WHEN s_4_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_4(51) WHEN s_4_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_4(52) WHEN s_4_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_4(53) WHEN s_4_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_4(54) WHEN s_4_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_4(55) WHEN s_4_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_4(56) WHEN s_4_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_4(57) WHEN s_4_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_4(58) WHEN s_4_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_4(59) WHEN s_4_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_4(60) WHEN s_4_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_4(61) WHEN s_4_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_4(62) WHEN s_4_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_4(63) WHEN s_4_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_4(64) WHEN s_4_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_4(65) WHEN s_4_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_4(66) WHEN s_4_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_4(67) WHEN s_4_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_4(68) WHEN s_4_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_4(69) WHEN s_4_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_4(70) WHEN s_4_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_4(71) WHEN s_4_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_4(72) WHEN s_4_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_4(73) WHEN s_4_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_4(74) WHEN s_4_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_4(75) WHEN s_4_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_4(76) WHEN s_4_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_4(77) WHEN s_4_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_4(78) WHEN s_4_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_4(79) WHEN s_4_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_4(80) WHEN s_4_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_4(81) WHEN s_4_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_4(82) WHEN s_4_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_4(83) WHEN s_4_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_4(84) WHEN s_4_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_4(85) WHEN s_4_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_4(86) WHEN s_4_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_4(87) WHEN s_4_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_4(88) WHEN s_4_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_4(89) WHEN s_4_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_4(90) WHEN s_4_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_4(91) WHEN s_4_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_4(92) WHEN s_4_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_4(93) WHEN s_4_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_4(94) WHEN s_4_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_4(95) WHEN s_4_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_4(96) WHEN s_4_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_4(97) WHEN s_4_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_4(98) WHEN s_4_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_4(99) WHEN s_4_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_4(100) WHEN s_4_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_4(101) WHEN s_4_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_4(102) WHEN s_4_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_4(103) WHEN s_4_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_4(104) WHEN s_4_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_4(105) WHEN s_4_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_4(106) WHEN s_4_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_4(107) WHEN s_4_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_4(108) WHEN s_4_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_4(109) WHEN s_4_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_4(110) WHEN s_4_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_4(111) WHEN s_4_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_4(112) WHEN s_4_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_4(113) WHEN s_4_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_4(114) WHEN s_4_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_4(115) WHEN s_4_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_4(116) WHEN s_4_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_4(117) WHEN s_4_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_4(118) WHEN s_4_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_4(119) WHEN s_4_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_4(120) WHEN s_4_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_4(121) WHEN s_4_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_4(122) WHEN s_4_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_4(123) WHEN s_4_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_4(124) WHEN s_4_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_4(125) WHEN s_4_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_4(126) WHEN s_4_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_4(127) WHEN s_4_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_4(128) WHEN s_4_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_4(129) WHEN s_4_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_4(130) WHEN s_4_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_4(131) WHEN s_4_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_4(132) WHEN s_4_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_4(133) WHEN s_4_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_4(134) WHEN s_4_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_4(135) WHEN s_4_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_4(136) WHEN s_4_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_4(137) WHEN s_4_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_4(138) WHEN s_4_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_4(139) WHEN s_4_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_4(140) WHEN s_4_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_4(141) WHEN s_4_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_4(142) WHEN s_4_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_4(143) WHEN s_4_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_4(144) WHEN s_4_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_4(145) WHEN s_4_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_4(146) WHEN s_4_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_4(147) WHEN s_4_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_4(148) WHEN s_4_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_4(149) WHEN s_4_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_4(150) WHEN s_4_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_4(151) WHEN s_4_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_4(152) WHEN s_4_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_4(153) WHEN s_4_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_4(154) WHEN s_4_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_4(155) WHEN s_4_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_4(156) WHEN s_4_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_4(157) WHEN s_4_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_4(158) WHEN s_4_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_4(159) WHEN s_4_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_4(160) WHEN s_4_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_4(161) WHEN s_4_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_4(162) WHEN s_4_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_4(163) WHEN s_4_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_4(164) WHEN s_4_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_4(165) WHEN s_4_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_4(166) WHEN s_4_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_4(167) WHEN s_4_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_4(168) WHEN s_4_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_4(169) WHEN s_4_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_4(170) WHEN s_4_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_4(171) WHEN s_4_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_4(172) WHEN s_4_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_4(173) WHEN s_4_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_4(174) WHEN s_4_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_4(175) WHEN s_4_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_4(176) WHEN s_4_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_4(177) WHEN s_4_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_4(178) WHEN s_4_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_4(179) WHEN s_4_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_4(180) WHEN s_4_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_4(181) WHEN s_4_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_4(182) WHEN s_4_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_4(183) WHEN s_4_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_4(184) WHEN s_4_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_4(185) WHEN s_4_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_4(186) WHEN s_4_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_4(187) WHEN s_4_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_4(188) WHEN s_4_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_4(189) WHEN s_4_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_4(190) WHEN s_4_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_4(191) WHEN s_4_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_4(192) WHEN s_4_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_4(193) WHEN s_4_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_4(194) WHEN s_4_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_4(195) WHEN s_4_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_4(196) WHEN s_4_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_4(197) WHEN s_4_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_4(198) WHEN s_4_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_4(199) WHEN s_4_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_4(200) WHEN s_4_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_4(201) WHEN s_4_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_4(202) WHEN s_4_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_4(203) WHEN s_4_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_4(204) WHEN s_4_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_4(205) WHEN s_4_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_4(206) WHEN s_4_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_4(207) WHEN s_4_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_4(208) WHEN s_4_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_4(209) WHEN s_4_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_4(210) WHEN s_4_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_4(211) WHEN s_4_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_4(212) WHEN s_4_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_4(213) WHEN s_4_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_4(214) WHEN s_4_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_4(215) WHEN s_4_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_4(216) WHEN s_4_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_4(217) WHEN s_4_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_4(218) WHEN s_4_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_4(219) WHEN s_4_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_4(220) WHEN s_4_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_4(221) WHEN s_4_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_4(222) WHEN s_4_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_4(223) WHEN s_4_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_4(224) WHEN s_4_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_4(225) WHEN s_4_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_4(226) WHEN s_4_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_4(227) WHEN s_4_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_4(228) WHEN s_4_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_4(229) WHEN s_4_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_4(230) WHEN s_4_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_4(231) WHEN s_4_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_4(232) WHEN s_4_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_4(233) WHEN s_4_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_4(234) WHEN s_4_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_4(235) WHEN s_4_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_4(236) WHEN s_4_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_4(237) WHEN s_4_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_4(238) WHEN s_4_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_4(239) WHEN s_4_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_4(240) WHEN s_4_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_4(241) WHEN s_4_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_4(242) WHEN s_4_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_4(243) WHEN s_4_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_4(244) WHEN s_4_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_4(245) WHEN s_4_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_4(246) WHEN s_4_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_4(247) WHEN s_4_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_4(248) WHEN s_4_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_4(249) WHEN s_4_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_4(250) WHEN s_4_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_4(251) WHEN s_4_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_4(252) WHEN s_4_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_4(253) WHEN s_4_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_4(254) WHEN s_4_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_4(255);

  out0_173 <= out0_172 XOR out0_171;

  b1_2 <= out0_173 XOR s_6_1;

  out0_174 <= b1_2 XOR s_7_1;

  
  out0_175 <= gmul2_3(0) WHEN s_3_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_3(1) WHEN s_3_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_3(2) WHEN s_3_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_3(3) WHEN s_3_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_3(4) WHEN s_3_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_3(5) WHEN s_3_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_3(6) WHEN s_3_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_3(7) WHEN s_3_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_3(8) WHEN s_3_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_3(9) WHEN s_3_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_3(10) WHEN s_3_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_3(11) WHEN s_3_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_3(12) WHEN s_3_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_3(13) WHEN s_3_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_3(14) WHEN s_3_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_3(15) WHEN s_3_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_3(16) WHEN s_3_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_3(17) WHEN s_3_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_3(18) WHEN s_3_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_3(19) WHEN s_3_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_3(20) WHEN s_3_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_3(21) WHEN s_3_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_3(22) WHEN s_3_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_3(23) WHEN s_3_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_3(24) WHEN s_3_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_3(25) WHEN s_3_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_3(26) WHEN s_3_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_3(27) WHEN s_3_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_3(28) WHEN s_3_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_3(29) WHEN s_3_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_3(30) WHEN s_3_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_3(31) WHEN s_3_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_3(32) WHEN s_3_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_3(33) WHEN s_3_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_3(34) WHEN s_3_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_3(35) WHEN s_3_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_3(36) WHEN s_3_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_3(37) WHEN s_3_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_3(38) WHEN s_3_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_3(39) WHEN s_3_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_3(40) WHEN s_3_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_3(41) WHEN s_3_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_3(42) WHEN s_3_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_3(43) WHEN s_3_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_3(44) WHEN s_3_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_3(45) WHEN s_3_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_3(46) WHEN s_3_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_3(47) WHEN s_3_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_3(48) WHEN s_3_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_3(49) WHEN s_3_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_3(50) WHEN s_3_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_3(51) WHEN s_3_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_3(52) WHEN s_3_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_3(53) WHEN s_3_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_3(54) WHEN s_3_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_3(55) WHEN s_3_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_3(56) WHEN s_3_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_3(57) WHEN s_3_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_3(58) WHEN s_3_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_3(59) WHEN s_3_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_3(60) WHEN s_3_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_3(61) WHEN s_3_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_3(62) WHEN s_3_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_3(63) WHEN s_3_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_3(64) WHEN s_3_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_3(65) WHEN s_3_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_3(66) WHEN s_3_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_3(67) WHEN s_3_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_3(68) WHEN s_3_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_3(69) WHEN s_3_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_3(70) WHEN s_3_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_3(71) WHEN s_3_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_3(72) WHEN s_3_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_3(73) WHEN s_3_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_3(74) WHEN s_3_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_3(75) WHEN s_3_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_3(76) WHEN s_3_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_3(77) WHEN s_3_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_3(78) WHEN s_3_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_3(79) WHEN s_3_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_3(80) WHEN s_3_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_3(81) WHEN s_3_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_3(82) WHEN s_3_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_3(83) WHEN s_3_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_3(84) WHEN s_3_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_3(85) WHEN s_3_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_3(86) WHEN s_3_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_3(87) WHEN s_3_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_3(88) WHEN s_3_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_3(89) WHEN s_3_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_3(90) WHEN s_3_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_3(91) WHEN s_3_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_3(92) WHEN s_3_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_3(93) WHEN s_3_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_3(94) WHEN s_3_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_3(95) WHEN s_3_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_3(96) WHEN s_3_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_3(97) WHEN s_3_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_3(98) WHEN s_3_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_3(99) WHEN s_3_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_3(100) WHEN s_3_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_3(101) WHEN s_3_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_3(102) WHEN s_3_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_3(103) WHEN s_3_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_3(104) WHEN s_3_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_3(105) WHEN s_3_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_3(106) WHEN s_3_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_3(107) WHEN s_3_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_3(108) WHEN s_3_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_3(109) WHEN s_3_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_3(110) WHEN s_3_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_3(111) WHEN s_3_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_3(112) WHEN s_3_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_3(113) WHEN s_3_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_3(114) WHEN s_3_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_3(115) WHEN s_3_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_3(116) WHEN s_3_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_3(117) WHEN s_3_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_3(118) WHEN s_3_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_3(119) WHEN s_3_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_3(120) WHEN s_3_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_3(121) WHEN s_3_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_3(122) WHEN s_3_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_3(123) WHEN s_3_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_3(124) WHEN s_3_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_3(125) WHEN s_3_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_3(126) WHEN s_3_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_3(127) WHEN s_3_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_3(128) WHEN s_3_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_3(129) WHEN s_3_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_3(130) WHEN s_3_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_3(131) WHEN s_3_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_3(132) WHEN s_3_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_3(133) WHEN s_3_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_3(134) WHEN s_3_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_3(135) WHEN s_3_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_3(136) WHEN s_3_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_3(137) WHEN s_3_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_3(138) WHEN s_3_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_3(139) WHEN s_3_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_3(140) WHEN s_3_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_3(141) WHEN s_3_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_3(142) WHEN s_3_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_3(143) WHEN s_3_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_3(144) WHEN s_3_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_3(145) WHEN s_3_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_3(146) WHEN s_3_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_3(147) WHEN s_3_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_3(148) WHEN s_3_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_3(149) WHEN s_3_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_3(150) WHEN s_3_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_3(151) WHEN s_3_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_3(152) WHEN s_3_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_3(153) WHEN s_3_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_3(154) WHEN s_3_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_3(155) WHEN s_3_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_3(156) WHEN s_3_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_3(157) WHEN s_3_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_3(158) WHEN s_3_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_3(159) WHEN s_3_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_3(160) WHEN s_3_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_3(161) WHEN s_3_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_3(162) WHEN s_3_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_3(163) WHEN s_3_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_3(164) WHEN s_3_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_3(165) WHEN s_3_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_3(166) WHEN s_3_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_3(167) WHEN s_3_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_3(168) WHEN s_3_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_3(169) WHEN s_3_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_3(170) WHEN s_3_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_3(171) WHEN s_3_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_3(172) WHEN s_3_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_3(173) WHEN s_3_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_3(174) WHEN s_3_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_3(175) WHEN s_3_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_3(176) WHEN s_3_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_3(177) WHEN s_3_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_3(178) WHEN s_3_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_3(179) WHEN s_3_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_3(180) WHEN s_3_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_3(181) WHEN s_3_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_3(182) WHEN s_3_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_3(183) WHEN s_3_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_3(184) WHEN s_3_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_3(185) WHEN s_3_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_3(186) WHEN s_3_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_3(187) WHEN s_3_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_3(188) WHEN s_3_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_3(189) WHEN s_3_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_3(190) WHEN s_3_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_3(191) WHEN s_3_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_3(192) WHEN s_3_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_3(193) WHEN s_3_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_3(194) WHEN s_3_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_3(195) WHEN s_3_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_3(196) WHEN s_3_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_3(197) WHEN s_3_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_3(198) WHEN s_3_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_3(199) WHEN s_3_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_3(200) WHEN s_3_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_3(201) WHEN s_3_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_3(202) WHEN s_3_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_3(203) WHEN s_3_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_3(204) WHEN s_3_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_3(205) WHEN s_3_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_3(206) WHEN s_3_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_3(207) WHEN s_3_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_3(208) WHEN s_3_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_3(209) WHEN s_3_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_3(210) WHEN s_3_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_3(211) WHEN s_3_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_3(212) WHEN s_3_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_3(213) WHEN s_3_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_3(214) WHEN s_3_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_3(215) WHEN s_3_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_3(216) WHEN s_3_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_3(217) WHEN s_3_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_3(218) WHEN s_3_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_3(219) WHEN s_3_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_3(220) WHEN s_3_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_3(221) WHEN s_3_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_3(222) WHEN s_3_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_3(223) WHEN s_3_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_3(224) WHEN s_3_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_3(225) WHEN s_3_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_3(226) WHEN s_3_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_3(227) WHEN s_3_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_3(228) WHEN s_3_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_3(229) WHEN s_3_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_3(230) WHEN s_3_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_3(231) WHEN s_3_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_3(232) WHEN s_3_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_3(233) WHEN s_3_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_3(234) WHEN s_3_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_3(235) WHEN s_3_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_3(236) WHEN s_3_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_3(237) WHEN s_3_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_3(238) WHEN s_3_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_3(239) WHEN s_3_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_3(240) WHEN s_3_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_3(241) WHEN s_3_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_3(242) WHEN s_3_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_3(243) WHEN s_3_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_3(244) WHEN s_3_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_3(245) WHEN s_3_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_3(246) WHEN s_3_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_3(247) WHEN s_3_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_3(248) WHEN s_3_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_3(249) WHEN s_3_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_3(250) WHEN s_3_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_3(251) WHEN s_3_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_3(252) WHEN s_3_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_3(253) WHEN s_3_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_3(254) WHEN s_3_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_3(255);

  
  out0_176 <= gmul3_3(0) WHEN s_0_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_3(1) WHEN s_0_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_3(2) WHEN s_0_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_3(3) WHEN s_0_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_3(4) WHEN s_0_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_3(5) WHEN s_0_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_3(6) WHEN s_0_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_3(7) WHEN s_0_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_3(8) WHEN s_0_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_3(9) WHEN s_0_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_3(10) WHEN s_0_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_3(11) WHEN s_0_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_3(12) WHEN s_0_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_3(13) WHEN s_0_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_3(14) WHEN s_0_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_3(15) WHEN s_0_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_3(16) WHEN s_0_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_3(17) WHEN s_0_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_3(18) WHEN s_0_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_3(19) WHEN s_0_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_3(20) WHEN s_0_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_3(21) WHEN s_0_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_3(22) WHEN s_0_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_3(23) WHEN s_0_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_3(24) WHEN s_0_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_3(25) WHEN s_0_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_3(26) WHEN s_0_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_3(27) WHEN s_0_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_3(28) WHEN s_0_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_3(29) WHEN s_0_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_3(30) WHEN s_0_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_3(31) WHEN s_0_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_3(32) WHEN s_0_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_3(33) WHEN s_0_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_3(34) WHEN s_0_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_3(35) WHEN s_0_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_3(36) WHEN s_0_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_3(37) WHEN s_0_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_3(38) WHEN s_0_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_3(39) WHEN s_0_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_3(40) WHEN s_0_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_3(41) WHEN s_0_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_3(42) WHEN s_0_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_3(43) WHEN s_0_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_3(44) WHEN s_0_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_3(45) WHEN s_0_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_3(46) WHEN s_0_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_3(47) WHEN s_0_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_3(48) WHEN s_0_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_3(49) WHEN s_0_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_3(50) WHEN s_0_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_3(51) WHEN s_0_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_3(52) WHEN s_0_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_3(53) WHEN s_0_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_3(54) WHEN s_0_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_3(55) WHEN s_0_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_3(56) WHEN s_0_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_3(57) WHEN s_0_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_3(58) WHEN s_0_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_3(59) WHEN s_0_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_3(60) WHEN s_0_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_3(61) WHEN s_0_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_3(62) WHEN s_0_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_3(63) WHEN s_0_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_3(64) WHEN s_0_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_3(65) WHEN s_0_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_3(66) WHEN s_0_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_3(67) WHEN s_0_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_3(68) WHEN s_0_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_3(69) WHEN s_0_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_3(70) WHEN s_0_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_3(71) WHEN s_0_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_3(72) WHEN s_0_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_3(73) WHEN s_0_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_3(74) WHEN s_0_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_3(75) WHEN s_0_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_3(76) WHEN s_0_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_3(77) WHEN s_0_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_3(78) WHEN s_0_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_3(79) WHEN s_0_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_3(80) WHEN s_0_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_3(81) WHEN s_0_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_3(82) WHEN s_0_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_3(83) WHEN s_0_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_3(84) WHEN s_0_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_3(85) WHEN s_0_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_3(86) WHEN s_0_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_3(87) WHEN s_0_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_3(88) WHEN s_0_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_3(89) WHEN s_0_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_3(90) WHEN s_0_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_3(91) WHEN s_0_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_3(92) WHEN s_0_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_3(93) WHEN s_0_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_3(94) WHEN s_0_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_3(95) WHEN s_0_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_3(96) WHEN s_0_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_3(97) WHEN s_0_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_3(98) WHEN s_0_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_3(99) WHEN s_0_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_3(100) WHEN s_0_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_3(101) WHEN s_0_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_3(102) WHEN s_0_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_3(103) WHEN s_0_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_3(104) WHEN s_0_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_3(105) WHEN s_0_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_3(106) WHEN s_0_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_3(107) WHEN s_0_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_3(108) WHEN s_0_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_3(109) WHEN s_0_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_3(110) WHEN s_0_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_3(111) WHEN s_0_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_3(112) WHEN s_0_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_3(113) WHEN s_0_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_3(114) WHEN s_0_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_3(115) WHEN s_0_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_3(116) WHEN s_0_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_3(117) WHEN s_0_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_3(118) WHEN s_0_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_3(119) WHEN s_0_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_3(120) WHEN s_0_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_3(121) WHEN s_0_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_3(122) WHEN s_0_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_3(123) WHEN s_0_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_3(124) WHEN s_0_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_3(125) WHEN s_0_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_3(126) WHEN s_0_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_3(127) WHEN s_0_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_3(128) WHEN s_0_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_3(129) WHEN s_0_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_3(130) WHEN s_0_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_3(131) WHEN s_0_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_3(132) WHEN s_0_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_3(133) WHEN s_0_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_3(134) WHEN s_0_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_3(135) WHEN s_0_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_3(136) WHEN s_0_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_3(137) WHEN s_0_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_3(138) WHEN s_0_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_3(139) WHEN s_0_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_3(140) WHEN s_0_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_3(141) WHEN s_0_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_3(142) WHEN s_0_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_3(143) WHEN s_0_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_3(144) WHEN s_0_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_3(145) WHEN s_0_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_3(146) WHEN s_0_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_3(147) WHEN s_0_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_3(148) WHEN s_0_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_3(149) WHEN s_0_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_3(150) WHEN s_0_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_3(151) WHEN s_0_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_3(152) WHEN s_0_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_3(153) WHEN s_0_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_3(154) WHEN s_0_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_3(155) WHEN s_0_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_3(156) WHEN s_0_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_3(157) WHEN s_0_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_3(158) WHEN s_0_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_3(159) WHEN s_0_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_3(160) WHEN s_0_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_3(161) WHEN s_0_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_3(162) WHEN s_0_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_3(163) WHEN s_0_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_3(164) WHEN s_0_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_3(165) WHEN s_0_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_3(166) WHEN s_0_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_3(167) WHEN s_0_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_3(168) WHEN s_0_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_3(169) WHEN s_0_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_3(170) WHEN s_0_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_3(171) WHEN s_0_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_3(172) WHEN s_0_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_3(173) WHEN s_0_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_3(174) WHEN s_0_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_3(175) WHEN s_0_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_3(176) WHEN s_0_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_3(177) WHEN s_0_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_3(178) WHEN s_0_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_3(179) WHEN s_0_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_3(180) WHEN s_0_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_3(181) WHEN s_0_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_3(182) WHEN s_0_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_3(183) WHEN s_0_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_3(184) WHEN s_0_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_3(185) WHEN s_0_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_3(186) WHEN s_0_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_3(187) WHEN s_0_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_3(188) WHEN s_0_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_3(189) WHEN s_0_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_3(190) WHEN s_0_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_3(191) WHEN s_0_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_3(192) WHEN s_0_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_3(193) WHEN s_0_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_3(194) WHEN s_0_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_3(195) WHEN s_0_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_3(196) WHEN s_0_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_3(197) WHEN s_0_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_3(198) WHEN s_0_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_3(199) WHEN s_0_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_3(200) WHEN s_0_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_3(201) WHEN s_0_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_3(202) WHEN s_0_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_3(203) WHEN s_0_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_3(204) WHEN s_0_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_3(205) WHEN s_0_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_3(206) WHEN s_0_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_3(207) WHEN s_0_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_3(208) WHEN s_0_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_3(209) WHEN s_0_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_3(210) WHEN s_0_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_3(211) WHEN s_0_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_3(212) WHEN s_0_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_3(213) WHEN s_0_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_3(214) WHEN s_0_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_3(215) WHEN s_0_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_3(216) WHEN s_0_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_3(217) WHEN s_0_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_3(218) WHEN s_0_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_3(219) WHEN s_0_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_3(220) WHEN s_0_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_3(221) WHEN s_0_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_3(222) WHEN s_0_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_3(223) WHEN s_0_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_3(224) WHEN s_0_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_3(225) WHEN s_0_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_3(226) WHEN s_0_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_3(227) WHEN s_0_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_3(228) WHEN s_0_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_3(229) WHEN s_0_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_3(230) WHEN s_0_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_3(231) WHEN s_0_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_3(232) WHEN s_0_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_3(233) WHEN s_0_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_3(234) WHEN s_0_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_3(235) WHEN s_0_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_3(236) WHEN s_0_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_3(237) WHEN s_0_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_3(238) WHEN s_0_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_3(239) WHEN s_0_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_3(240) WHEN s_0_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_3(241) WHEN s_0_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_3(242) WHEN s_0_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_3(243) WHEN s_0_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_3(244) WHEN s_0_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_3(245) WHEN s_0_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_3(246) WHEN s_0_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_3(247) WHEN s_0_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_3(248) WHEN s_0_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_3(249) WHEN s_0_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_3(250) WHEN s_0_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_3(251) WHEN s_0_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_3(252) WHEN s_0_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_3(253) WHEN s_0_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_3(254) WHEN s_0_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_3(255);

  out0_177 <= out0_176 XOR s_1_1;

  b4_3 <= out0_177 XOR s_2_1;

  out0_178 <= b4_3 XOR out0_175;

  
  out0_179 <= gmul3_2(0) WHEN s_3_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_2(1) WHEN s_3_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_2(2) WHEN s_3_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_2(3) WHEN s_3_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_2(4) WHEN s_3_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_2(5) WHEN s_3_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_2(6) WHEN s_3_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_2(7) WHEN s_3_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_2(8) WHEN s_3_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_2(9) WHEN s_3_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_2(10) WHEN s_3_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_2(11) WHEN s_3_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_2(12) WHEN s_3_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_2(13) WHEN s_3_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_2(14) WHEN s_3_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_2(15) WHEN s_3_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_2(16) WHEN s_3_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_2(17) WHEN s_3_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_2(18) WHEN s_3_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_2(19) WHEN s_3_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_2(20) WHEN s_3_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_2(21) WHEN s_3_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_2(22) WHEN s_3_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_2(23) WHEN s_3_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_2(24) WHEN s_3_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_2(25) WHEN s_3_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_2(26) WHEN s_3_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_2(27) WHEN s_3_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_2(28) WHEN s_3_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_2(29) WHEN s_3_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_2(30) WHEN s_3_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_2(31) WHEN s_3_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_2(32) WHEN s_3_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_2(33) WHEN s_3_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_2(34) WHEN s_3_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_2(35) WHEN s_3_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_2(36) WHEN s_3_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_2(37) WHEN s_3_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_2(38) WHEN s_3_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_2(39) WHEN s_3_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_2(40) WHEN s_3_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_2(41) WHEN s_3_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_2(42) WHEN s_3_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_2(43) WHEN s_3_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_2(44) WHEN s_3_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_2(45) WHEN s_3_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_2(46) WHEN s_3_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_2(47) WHEN s_3_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_2(48) WHEN s_3_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_2(49) WHEN s_3_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_2(50) WHEN s_3_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_2(51) WHEN s_3_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_2(52) WHEN s_3_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_2(53) WHEN s_3_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_2(54) WHEN s_3_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_2(55) WHEN s_3_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_2(56) WHEN s_3_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_2(57) WHEN s_3_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_2(58) WHEN s_3_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_2(59) WHEN s_3_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_2(60) WHEN s_3_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_2(61) WHEN s_3_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_2(62) WHEN s_3_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_2(63) WHEN s_3_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_2(64) WHEN s_3_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_2(65) WHEN s_3_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_2(66) WHEN s_3_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_2(67) WHEN s_3_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_2(68) WHEN s_3_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_2(69) WHEN s_3_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_2(70) WHEN s_3_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_2(71) WHEN s_3_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_2(72) WHEN s_3_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_2(73) WHEN s_3_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_2(74) WHEN s_3_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_2(75) WHEN s_3_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_2(76) WHEN s_3_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_2(77) WHEN s_3_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_2(78) WHEN s_3_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_2(79) WHEN s_3_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_2(80) WHEN s_3_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_2(81) WHEN s_3_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_2(82) WHEN s_3_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_2(83) WHEN s_3_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_2(84) WHEN s_3_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_2(85) WHEN s_3_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_2(86) WHEN s_3_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_2(87) WHEN s_3_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_2(88) WHEN s_3_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_2(89) WHEN s_3_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_2(90) WHEN s_3_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_2(91) WHEN s_3_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_2(92) WHEN s_3_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_2(93) WHEN s_3_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_2(94) WHEN s_3_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_2(95) WHEN s_3_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_2(96) WHEN s_3_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_2(97) WHEN s_3_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_2(98) WHEN s_3_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_2(99) WHEN s_3_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_2(100) WHEN s_3_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_2(101) WHEN s_3_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_2(102) WHEN s_3_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_2(103) WHEN s_3_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_2(104) WHEN s_3_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_2(105) WHEN s_3_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_2(106) WHEN s_3_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_2(107) WHEN s_3_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_2(108) WHEN s_3_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_2(109) WHEN s_3_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_2(110) WHEN s_3_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_2(111) WHEN s_3_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_2(112) WHEN s_3_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_2(113) WHEN s_3_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_2(114) WHEN s_3_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_2(115) WHEN s_3_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_2(116) WHEN s_3_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_2(117) WHEN s_3_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_2(118) WHEN s_3_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_2(119) WHEN s_3_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_2(120) WHEN s_3_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_2(121) WHEN s_3_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_2(122) WHEN s_3_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_2(123) WHEN s_3_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_2(124) WHEN s_3_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_2(125) WHEN s_3_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_2(126) WHEN s_3_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_2(127) WHEN s_3_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_2(128) WHEN s_3_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_2(129) WHEN s_3_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_2(130) WHEN s_3_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_2(131) WHEN s_3_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_2(132) WHEN s_3_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_2(133) WHEN s_3_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_2(134) WHEN s_3_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_2(135) WHEN s_3_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_2(136) WHEN s_3_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_2(137) WHEN s_3_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_2(138) WHEN s_3_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_2(139) WHEN s_3_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_2(140) WHEN s_3_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_2(141) WHEN s_3_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_2(142) WHEN s_3_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_2(143) WHEN s_3_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_2(144) WHEN s_3_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_2(145) WHEN s_3_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_2(146) WHEN s_3_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_2(147) WHEN s_3_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_2(148) WHEN s_3_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_2(149) WHEN s_3_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_2(150) WHEN s_3_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_2(151) WHEN s_3_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_2(152) WHEN s_3_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_2(153) WHEN s_3_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_2(154) WHEN s_3_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_2(155) WHEN s_3_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_2(156) WHEN s_3_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_2(157) WHEN s_3_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_2(158) WHEN s_3_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_2(159) WHEN s_3_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_2(160) WHEN s_3_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_2(161) WHEN s_3_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_2(162) WHEN s_3_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_2(163) WHEN s_3_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_2(164) WHEN s_3_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_2(165) WHEN s_3_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_2(166) WHEN s_3_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_2(167) WHEN s_3_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_2(168) WHEN s_3_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_2(169) WHEN s_3_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_2(170) WHEN s_3_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_2(171) WHEN s_3_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_2(172) WHEN s_3_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_2(173) WHEN s_3_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_2(174) WHEN s_3_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_2(175) WHEN s_3_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_2(176) WHEN s_3_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_2(177) WHEN s_3_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_2(178) WHEN s_3_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_2(179) WHEN s_3_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_2(180) WHEN s_3_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_2(181) WHEN s_3_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_2(182) WHEN s_3_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_2(183) WHEN s_3_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_2(184) WHEN s_3_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_2(185) WHEN s_3_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_2(186) WHEN s_3_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_2(187) WHEN s_3_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_2(188) WHEN s_3_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_2(189) WHEN s_3_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_2(190) WHEN s_3_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_2(191) WHEN s_3_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_2(192) WHEN s_3_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_2(193) WHEN s_3_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_2(194) WHEN s_3_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_2(195) WHEN s_3_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_2(196) WHEN s_3_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_2(197) WHEN s_3_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_2(198) WHEN s_3_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_2(199) WHEN s_3_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_2(200) WHEN s_3_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_2(201) WHEN s_3_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_2(202) WHEN s_3_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_2(203) WHEN s_3_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_2(204) WHEN s_3_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_2(205) WHEN s_3_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_2(206) WHEN s_3_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_2(207) WHEN s_3_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_2(208) WHEN s_3_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_2(209) WHEN s_3_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_2(210) WHEN s_3_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_2(211) WHEN s_3_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_2(212) WHEN s_3_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_2(213) WHEN s_3_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_2(214) WHEN s_3_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_2(215) WHEN s_3_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_2(216) WHEN s_3_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_2(217) WHEN s_3_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_2(218) WHEN s_3_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_2(219) WHEN s_3_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_2(220) WHEN s_3_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_2(221) WHEN s_3_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_2(222) WHEN s_3_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_2(223) WHEN s_3_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_2(224) WHEN s_3_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_2(225) WHEN s_3_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_2(226) WHEN s_3_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_2(227) WHEN s_3_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_2(228) WHEN s_3_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_2(229) WHEN s_3_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_2(230) WHEN s_3_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_2(231) WHEN s_3_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_2(232) WHEN s_3_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_2(233) WHEN s_3_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_2(234) WHEN s_3_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_2(235) WHEN s_3_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_2(236) WHEN s_3_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_2(237) WHEN s_3_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_2(238) WHEN s_3_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_2(239) WHEN s_3_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_2(240) WHEN s_3_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_2(241) WHEN s_3_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_2(242) WHEN s_3_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_2(243) WHEN s_3_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_2(244) WHEN s_3_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_2(245) WHEN s_3_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_2(246) WHEN s_3_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_2(247) WHEN s_3_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_2(248) WHEN s_3_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_2(249) WHEN s_3_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_2(250) WHEN s_3_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_2(251) WHEN s_3_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_2(252) WHEN s_3_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_2(253) WHEN s_3_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_2(254) WHEN s_3_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_2(255);

  
  out0_180 <= gmul2_2(0) WHEN s_2_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_2(1) WHEN s_2_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_2(2) WHEN s_2_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_2(3) WHEN s_2_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_2(4) WHEN s_2_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_2(5) WHEN s_2_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_2(6) WHEN s_2_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_2(7) WHEN s_2_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_2(8) WHEN s_2_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_2(9) WHEN s_2_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_2(10) WHEN s_2_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_2(11) WHEN s_2_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_2(12) WHEN s_2_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_2(13) WHEN s_2_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_2(14) WHEN s_2_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_2(15) WHEN s_2_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_2(16) WHEN s_2_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_2(17) WHEN s_2_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_2(18) WHEN s_2_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_2(19) WHEN s_2_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_2(20) WHEN s_2_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_2(21) WHEN s_2_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_2(22) WHEN s_2_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_2(23) WHEN s_2_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_2(24) WHEN s_2_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_2(25) WHEN s_2_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_2(26) WHEN s_2_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_2(27) WHEN s_2_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_2(28) WHEN s_2_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_2(29) WHEN s_2_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_2(30) WHEN s_2_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_2(31) WHEN s_2_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_2(32) WHEN s_2_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_2(33) WHEN s_2_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_2(34) WHEN s_2_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_2(35) WHEN s_2_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_2(36) WHEN s_2_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_2(37) WHEN s_2_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_2(38) WHEN s_2_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_2(39) WHEN s_2_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_2(40) WHEN s_2_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_2(41) WHEN s_2_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_2(42) WHEN s_2_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_2(43) WHEN s_2_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_2(44) WHEN s_2_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_2(45) WHEN s_2_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_2(46) WHEN s_2_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_2(47) WHEN s_2_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_2(48) WHEN s_2_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_2(49) WHEN s_2_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_2(50) WHEN s_2_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_2(51) WHEN s_2_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_2(52) WHEN s_2_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_2(53) WHEN s_2_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_2(54) WHEN s_2_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_2(55) WHEN s_2_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_2(56) WHEN s_2_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_2(57) WHEN s_2_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_2(58) WHEN s_2_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_2(59) WHEN s_2_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_2(60) WHEN s_2_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_2(61) WHEN s_2_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_2(62) WHEN s_2_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_2(63) WHEN s_2_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_2(64) WHEN s_2_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_2(65) WHEN s_2_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_2(66) WHEN s_2_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_2(67) WHEN s_2_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_2(68) WHEN s_2_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_2(69) WHEN s_2_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_2(70) WHEN s_2_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_2(71) WHEN s_2_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_2(72) WHEN s_2_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_2(73) WHEN s_2_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_2(74) WHEN s_2_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_2(75) WHEN s_2_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_2(76) WHEN s_2_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_2(77) WHEN s_2_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_2(78) WHEN s_2_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_2(79) WHEN s_2_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_2(80) WHEN s_2_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_2(81) WHEN s_2_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_2(82) WHEN s_2_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_2(83) WHEN s_2_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_2(84) WHEN s_2_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_2(85) WHEN s_2_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_2(86) WHEN s_2_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_2(87) WHEN s_2_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_2(88) WHEN s_2_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_2(89) WHEN s_2_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_2(90) WHEN s_2_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_2(91) WHEN s_2_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_2(92) WHEN s_2_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_2(93) WHEN s_2_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_2(94) WHEN s_2_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_2(95) WHEN s_2_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_2(96) WHEN s_2_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_2(97) WHEN s_2_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_2(98) WHEN s_2_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_2(99) WHEN s_2_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_2(100) WHEN s_2_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_2(101) WHEN s_2_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_2(102) WHEN s_2_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_2(103) WHEN s_2_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_2(104) WHEN s_2_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_2(105) WHEN s_2_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_2(106) WHEN s_2_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_2(107) WHEN s_2_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_2(108) WHEN s_2_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_2(109) WHEN s_2_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_2(110) WHEN s_2_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_2(111) WHEN s_2_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_2(112) WHEN s_2_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_2(113) WHEN s_2_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_2(114) WHEN s_2_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_2(115) WHEN s_2_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_2(116) WHEN s_2_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_2(117) WHEN s_2_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_2(118) WHEN s_2_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_2(119) WHEN s_2_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_2(120) WHEN s_2_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_2(121) WHEN s_2_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_2(122) WHEN s_2_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_2(123) WHEN s_2_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_2(124) WHEN s_2_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_2(125) WHEN s_2_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_2(126) WHEN s_2_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_2(127) WHEN s_2_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_2(128) WHEN s_2_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_2(129) WHEN s_2_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_2(130) WHEN s_2_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_2(131) WHEN s_2_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_2(132) WHEN s_2_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_2(133) WHEN s_2_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_2(134) WHEN s_2_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_2(135) WHEN s_2_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_2(136) WHEN s_2_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_2(137) WHEN s_2_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_2(138) WHEN s_2_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_2(139) WHEN s_2_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_2(140) WHEN s_2_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_2(141) WHEN s_2_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_2(142) WHEN s_2_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_2(143) WHEN s_2_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_2(144) WHEN s_2_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_2(145) WHEN s_2_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_2(146) WHEN s_2_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_2(147) WHEN s_2_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_2(148) WHEN s_2_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_2(149) WHEN s_2_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_2(150) WHEN s_2_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_2(151) WHEN s_2_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_2(152) WHEN s_2_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_2(153) WHEN s_2_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_2(154) WHEN s_2_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_2(155) WHEN s_2_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_2(156) WHEN s_2_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_2(157) WHEN s_2_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_2(158) WHEN s_2_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_2(159) WHEN s_2_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_2(160) WHEN s_2_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_2(161) WHEN s_2_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_2(162) WHEN s_2_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_2(163) WHEN s_2_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_2(164) WHEN s_2_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_2(165) WHEN s_2_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_2(166) WHEN s_2_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_2(167) WHEN s_2_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_2(168) WHEN s_2_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_2(169) WHEN s_2_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_2(170) WHEN s_2_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_2(171) WHEN s_2_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_2(172) WHEN s_2_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_2(173) WHEN s_2_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_2(174) WHEN s_2_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_2(175) WHEN s_2_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_2(176) WHEN s_2_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_2(177) WHEN s_2_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_2(178) WHEN s_2_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_2(179) WHEN s_2_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_2(180) WHEN s_2_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_2(181) WHEN s_2_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_2(182) WHEN s_2_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_2(183) WHEN s_2_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_2(184) WHEN s_2_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_2(185) WHEN s_2_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_2(186) WHEN s_2_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_2(187) WHEN s_2_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_2(188) WHEN s_2_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_2(189) WHEN s_2_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_2(190) WHEN s_2_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_2(191) WHEN s_2_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_2(192) WHEN s_2_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_2(193) WHEN s_2_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_2(194) WHEN s_2_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_2(195) WHEN s_2_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_2(196) WHEN s_2_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_2(197) WHEN s_2_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_2(198) WHEN s_2_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_2(199) WHEN s_2_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_2(200) WHEN s_2_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_2(201) WHEN s_2_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_2(202) WHEN s_2_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_2(203) WHEN s_2_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_2(204) WHEN s_2_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_2(205) WHEN s_2_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_2(206) WHEN s_2_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_2(207) WHEN s_2_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_2(208) WHEN s_2_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_2(209) WHEN s_2_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_2(210) WHEN s_2_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_2(211) WHEN s_2_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_2(212) WHEN s_2_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_2(213) WHEN s_2_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_2(214) WHEN s_2_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_2(215) WHEN s_2_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_2(216) WHEN s_2_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_2(217) WHEN s_2_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_2(218) WHEN s_2_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_2(219) WHEN s_2_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_2(220) WHEN s_2_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_2(221) WHEN s_2_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_2(222) WHEN s_2_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_2(223) WHEN s_2_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_2(224) WHEN s_2_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_2(225) WHEN s_2_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_2(226) WHEN s_2_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_2(227) WHEN s_2_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_2(228) WHEN s_2_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_2(229) WHEN s_2_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_2(230) WHEN s_2_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_2(231) WHEN s_2_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_2(232) WHEN s_2_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_2(233) WHEN s_2_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_2(234) WHEN s_2_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_2(235) WHEN s_2_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_2(236) WHEN s_2_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_2(237) WHEN s_2_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_2(238) WHEN s_2_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_2(239) WHEN s_2_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_2(240) WHEN s_2_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_2(241) WHEN s_2_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_2(242) WHEN s_2_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_2(243) WHEN s_2_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_2(244) WHEN s_2_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_2(245) WHEN s_2_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_2(246) WHEN s_2_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_2(247) WHEN s_2_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_2(248) WHEN s_2_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_2(249) WHEN s_2_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_2(250) WHEN s_2_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_2(251) WHEN s_2_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_2(252) WHEN s_2_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_2(253) WHEN s_2_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_2(254) WHEN s_2_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_2(255);

  out0_181 <= s_0_1 XOR s_1_1;

  b3_3 <= out0_181 XOR out0_180;

  out0_182 <= b3_3 XOR out0_179;

  
  out0_183 <= gmul3_1(0) WHEN s_2_1 = to_unsigned(16#01#, 8) ELSE
      gmul3_1(1) WHEN s_2_1 = to_unsigned(16#02#, 8) ELSE
      gmul3_1(2) WHEN s_2_1 = to_unsigned(16#03#, 8) ELSE
      gmul3_1(3) WHEN s_2_1 = to_unsigned(16#04#, 8) ELSE
      gmul3_1(4) WHEN s_2_1 = to_unsigned(16#05#, 8) ELSE
      gmul3_1(5) WHEN s_2_1 = to_unsigned(16#06#, 8) ELSE
      gmul3_1(6) WHEN s_2_1 = to_unsigned(16#07#, 8) ELSE
      gmul3_1(7) WHEN s_2_1 = to_unsigned(16#08#, 8) ELSE
      gmul3_1(8) WHEN s_2_1 = to_unsigned(16#09#, 8) ELSE
      gmul3_1(9) WHEN s_2_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3_1(10) WHEN s_2_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3_1(11) WHEN s_2_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3_1(12) WHEN s_2_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3_1(13) WHEN s_2_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3_1(14) WHEN s_2_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3_1(15) WHEN s_2_1 = to_unsigned(16#10#, 8) ELSE
      gmul3_1(16) WHEN s_2_1 = to_unsigned(16#11#, 8) ELSE
      gmul3_1(17) WHEN s_2_1 = to_unsigned(16#12#, 8) ELSE
      gmul3_1(18) WHEN s_2_1 = to_unsigned(16#13#, 8) ELSE
      gmul3_1(19) WHEN s_2_1 = to_unsigned(16#14#, 8) ELSE
      gmul3_1(20) WHEN s_2_1 = to_unsigned(16#15#, 8) ELSE
      gmul3_1(21) WHEN s_2_1 = to_unsigned(16#16#, 8) ELSE
      gmul3_1(22) WHEN s_2_1 = to_unsigned(16#17#, 8) ELSE
      gmul3_1(23) WHEN s_2_1 = to_unsigned(16#18#, 8) ELSE
      gmul3_1(24) WHEN s_2_1 = to_unsigned(16#19#, 8) ELSE
      gmul3_1(25) WHEN s_2_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3_1(26) WHEN s_2_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3_1(27) WHEN s_2_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3_1(28) WHEN s_2_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3_1(29) WHEN s_2_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3_1(30) WHEN s_2_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3_1(31) WHEN s_2_1 = to_unsigned(16#20#, 8) ELSE
      gmul3_1(32) WHEN s_2_1 = to_unsigned(16#21#, 8) ELSE
      gmul3_1(33) WHEN s_2_1 = to_unsigned(16#22#, 8) ELSE
      gmul3_1(34) WHEN s_2_1 = to_unsigned(16#23#, 8) ELSE
      gmul3_1(35) WHEN s_2_1 = to_unsigned(16#24#, 8) ELSE
      gmul3_1(36) WHEN s_2_1 = to_unsigned(16#25#, 8) ELSE
      gmul3_1(37) WHEN s_2_1 = to_unsigned(16#26#, 8) ELSE
      gmul3_1(38) WHEN s_2_1 = to_unsigned(16#27#, 8) ELSE
      gmul3_1(39) WHEN s_2_1 = to_unsigned(16#28#, 8) ELSE
      gmul3_1(40) WHEN s_2_1 = to_unsigned(16#29#, 8) ELSE
      gmul3_1(41) WHEN s_2_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3_1(42) WHEN s_2_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3_1(43) WHEN s_2_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3_1(44) WHEN s_2_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3_1(45) WHEN s_2_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3_1(46) WHEN s_2_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3_1(47) WHEN s_2_1 = to_unsigned(16#30#, 8) ELSE
      gmul3_1(48) WHEN s_2_1 = to_unsigned(16#31#, 8) ELSE
      gmul3_1(49) WHEN s_2_1 = to_unsigned(16#32#, 8) ELSE
      gmul3_1(50) WHEN s_2_1 = to_unsigned(16#33#, 8) ELSE
      gmul3_1(51) WHEN s_2_1 = to_unsigned(16#34#, 8) ELSE
      gmul3_1(52) WHEN s_2_1 = to_unsigned(16#35#, 8) ELSE
      gmul3_1(53) WHEN s_2_1 = to_unsigned(16#36#, 8) ELSE
      gmul3_1(54) WHEN s_2_1 = to_unsigned(16#37#, 8) ELSE
      gmul3_1(55) WHEN s_2_1 = to_unsigned(16#38#, 8) ELSE
      gmul3_1(56) WHEN s_2_1 = to_unsigned(16#39#, 8) ELSE
      gmul3_1(57) WHEN s_2_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3_1(58) WHEN s_2_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3_1(59) WHEN s_2_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3_1(60) WHEN s_2_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3_1(61) WHEN s_2_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3_1(62) WHEN s_2_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3_1(63) WHEN s_2_1 = to_unsigned(16#40#, 8) ELSE
      gmul3_1(64) WHEN s_2_1 = to_unsigned(16#41#, 8) ELSE
      gmul3_1(65) WHEN s_2_1 = to_unsigned(16#42#, 8) ELSE
      gmul3_1(66) WHEN s_2_1 = to_unsigned(16#43#, 8) ELSE
      gmul3_1(67) WHEN s_2_1 = to_unsigned(16#44#, 8) ELSE
      gmul3_1(68) WHEN s_2_1 = to_unsigned(16#45#, 8) ELSE
      gmul3_1(69) WHEN s_2_1 = to_unsigned(16#46#, 8) ELSE
      gmul3_1(70) WHEN s_2_1 = to_unsigned(16#47#, 8) ELSE
      gmul3_1(71) WHEN s_2_1 = to_unsigned(16#48#, 8) ELSE
      gmul3_1(72) WHEN s_2_1 = to_unsigned(16#49#, 8) ELSE
      gmul3_1(73) WHEN s_2_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3_1(74) WHEN s_2_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3_1(75) WHEN s_2_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3_1(76) WHEN s_2_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3_1(77) WHEN s_2_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3_1(78) WHEN s_2_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3_1(79) WHEN s_2_1 = to_unsigned(16#50#, 8) ELSE
      gmul3_1(80) WHEN s_2_1 = to_unsigned(16#51#, 8) ELSE
      gmul3_1(81) WHEN s_2_1 = to_unsigned(16#52#, 8) ELSE
      gmul3_1(82) WHEN s_2_1 = to_unsigned(16#53#, 8) ELSE
      gmul3_1(83) WHEN s_2_1 = to_unsigned(16#54#, 8) ELSE
      gmul3_1(84) WHEN s_2_1 = to_unsigned(16#55#, 8) ELSE
      gmul3_1(85) WHEN s_2_1 = to_unsigned(16#56#, 8) ELSE
      gmul3_1(86) WHEN s_2_1 = to_unsigned(16#57#, 8) ELSE
      gmul3_1(87) WHEN s_2_1 = to_unsigned(16#58#, 8) ELSE
      gmul3_1(88) WHEN s_2_1 = to_unsigned(16#59#, 8) ELSE
      gmul3_1(89) WHEN s_2_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3_1(90) WHEN s_2_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3_1(91) WHEN s_2_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3_1(92) WHEN s_2_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3_1(93) WHEN s_2_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3_1(94) WHEN s_2_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3_1(95) WHEN s_2_1 = to_unsigned(16#60#, 8) ELSE
      gmul3_1(96) WHEN s_2_1 = to_unsigned(16#61#, 8) ELSE
      gmul3_1(97) WHEN s_2_1 = to_unsigned(16#62#, 8) ELSE
      gmul3_1(98) WHEN s_2_1 = to_unsigned(16#63#, 8) ELSE
      gmul3_1(99) WHEN s_2_1 = to_unsigned(16#64#, 8) ELSE
      gmul3_1(100) WHEN s_2_1 = to_unsigned(16#65#, 8) ELSE
      gmul3_1(101) WHEN s_2_1 = to_unsigned(16#66#, 8) ELSE
      gmul3_1(102) WHEN s_2_1 = to_unsigned(16#67#, 8) ELSE
      gmul3_1(103) WHEN s_2_1 = to_unsigned(16#68#, 8) ELSE
      gmul3_1(104) WHEN s_2_1 = to_unsigned(16#69#, 8) ELSE
      gmul3_1(105) WHEN s_2_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3_1(106) WHEN s_2_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3_1(107) WHEN s_2_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3_1(108) WHEN s_2_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3_1(109) WHEN s_2_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3_1(110) WHEN s_2_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3_1(111) WHEN s_2_1 = to_unsigned(16#70#, 8) ELSE
      gmul3_1(112) WHEN s_2_1 = to_unsigned(16#71#, 8) ELSE
      gmul3_1(113) WHEN s_2_1 = to_unsigned(16#72#, 8) ELSE
      gmul3_1(114) WHEN s_2_1 = to_unsigned(16#73#, 8) ELSE
      gmul3_1(115) WHEN s_2_1 = to_unsigned(16#74#, 8) ELSE
      gmul3_1(116) WHEN s_2_1 = to_unsigned(16#75#, 8) ELSE
      gmul3_1(117) WHEN s_2_1 = to_unsigned(16#76#, 8) ELSE
      gmul3_1(118) WHEN s_2_1 = to_unsigned(16#77#, 8) ELSE
      gmul3_1(119) WHEN s_2_1 = to_unsigned(16#78#, 8) ELSE
      gmul3_1(120) WHEN s_2_1 = to_unsigned(16#79#, 8) ELSE
      gmul3_1(121) WHEN s_2_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3_1(122) WHEN s_2_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3_1(123) WHEN s_2_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3_1(124) WHEN s_2_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3_1(125) WHEN s_2_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3_1(126) WHEN s_2_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3_1(127) WHEN s_2_1 = to_unsigned(16#80#, 8) ELSE
      gmul3_1(128) WHEN s_2_1 = to_unsigned(16#81#, 8) ELSE
      gmul3_1(129) WHEN s_2_1 = to_unsigned(16#82#, 8) ELSE
      gmul3_1(130) WHEN s_2_1 = to_unsigned(16#83#, 8) ELSE
      gmul3_1(131) WHEN s_2_1 = to_unsigned(16#84#, 8) ELSE
      gmul3_1(132) WHEN s_2_1 = to_unsigned(16#85#, 8) ELSE
      gmul3_1(133) WHEN s_2_1 = to_unsigned(16#86#, 8) ELSE
      gmul3_1(134) WHEN s_2_1 = to_unsigned(16#87#, 8) ELSE
      gmul3_1(135) WHEN s_2_1 = to_unsigned(16#88#, 8) ELSE
      gmul3_1(136) WHEN s_2_1 = to_unsigned(16#89#, 8) ELSE
      gmul3_1(137) WHEN s_2_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3_1(138) WHEN s_2_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3_1(139) WHEN s_2_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3_1(140) WHEN s_2_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3_1(141) WHEN s_2_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3_1(142) WHEN s_2_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3_1(143) WHEN s_2_1 = to_unsigned(16#90#, 8) ELSE
      gmul3_1(144) WHEN s_2_1 = to_unsigned(16#91#, 8) ELSE
      gmul3_1(145) WHEN s_2_1 = to_unsigned(16#92#, 8) ELSE
      gmul3_1(146) WHEN s_2_1 = to_unsigned(16#93#, 8) ELSE
      gmul3_1(147) WHEN s_2_1 = to_unsigned(16#94#, 8) ELSE
      gmul3_1(148) WHEN s_2_1 = to_unsigned(16#95#, 8) ELSE
      gmul3_1(149) WHEN s_2_1 = to_unsigned(16#96#, 8) ELSE
      gmul3_1(150) WHEN s_2_1 = to_unsigned(16#97#, 8) ELSE
      gmul3_1(151) WHEN s_2_1 = to_unsigned(16#98#, 8) ELSE
      gmul3_1(152) WHEN s_2_1 = to_unsigned(16#99#, 8) ELSE
      gmul3_1(153) WHEN s_2_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3_1(154) WHEN s_2_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3_1(155) WHEN s_2_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3_1(156) WHEN s_2_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3_1(157) WHEN s_2_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3_1(158) WHEN s_2_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3_1(159) WHEN s_2_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3_1(160) WHEN s_2_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3_1(161) WHEN s_2_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3_1(162) WHEN s_2_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3_1(163) WHEN s_2_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3_1(164) WHEN s_2_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3_1(165) WHEN s_2_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3_1(166) WHEN s_2_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3_1(167) WHEN s_2_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3_1(168) WHEN s_2_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3_1(169) WHEN s_2_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3_1(170) WHEN s_2_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3_1(171) WHEN s_2_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3_1(172) WHEN s_2_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3_1(173) WHEN s_2_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3_1(174) WHEN s_2_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3_1(175) WHEN s_2_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3_1(176) WHEN s_2_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3_1(177) WHEN s_2_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3_1(178) WHEN s_2_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3_1(179) WHEN s_2_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3_1(180) WHEN s_2_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3_1(181) WHEN s_2_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3_1(182) WHEN s_2_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3_1(183) WHEN s_2_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3_1(184) WHEN s_2_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3_1(185) WHEN s_2_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3_1(186) WHEN s_2_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3_1(187) WHEN s_2_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3_1(188) WHEN s_2_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3_1(189) WHEN s_2_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3_1(190) WHEN s_2_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3_1(191) WHEN s_2_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3_1(192) WHEN s_2_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3_1(193) WHEN s_2_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3_1(194) WHEN s_2_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3_1(195) WHEN s_2_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3_1(196) WHEN s_2_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3_1(197) WHEN s_2_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3_1(198) WHEN s_2_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3_1(199) WHEN s_2_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3_1(200) WHEN s_2_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3_1(201) WHEN s_2_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3_1(202) WHEN s_2_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3_1(203) WHEN s_2_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3_1(204) WHEN s_2_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3_1(205) WHEN s_2_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3_1(206) WHEN s_2_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3_1(207) WHEN s_2_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3_1(208) WHEN s_2_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3_1(209) WHEN s_2_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3_1(210) WHEN s_2_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3_1(211) WHEN s_2_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3_1(212) WHEN s_2_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3_1(213) WHEN s_2_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3_1(214) WHEN s_2_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3_1(215) WHEN s_2_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3_1(216) WHEN s_2_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3_1(217) WHEN s_2_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3_1(218) WHEN s_2_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3_1(219) WHEN s_2_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3_1(220) WHEN s_2_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3_1(221) WHEN s_2_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3_1(222) WHEN s_2_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3_1(223) WHEN s_2_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3_1(224) WHEN s_2_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3_1(225) WHEN s_2_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3_1(226) WHEN s_2_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3_1(227) WHEN s_2_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3_1(228) WHEN s_2_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3_1(229) WHEN s_2_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3_1(230) WHEN s_2_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3_1(231) WHEN s_2_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3_1(232) WHEN s_2_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3_1(233) WHEN s_2_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3_1(234) WHEN s_2_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3_1(235) WHEN s_2_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3_1(236) WHEN s_2_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3_1(237) WHEN s_2_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3_1(238) WHEN s_2_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3_1(239) WHEN s_2_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3_1(240) WHEN s_2_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3_1(241) WHEN s_2_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3_1(242) WHEN s_2_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3_1(243) WHEN s_2_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3_1(244) WHEN s_2_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3_1(245) WHEN s_2_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3_1(246) WHEN s_2_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3_1(247) WHEN s_2_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3_1(248) WHEN s_2_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3_1(249) WHEN s_2_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3_1(250) WHEN s_2_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3_1(251) WHEN s_2_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3_1(252) WHEN s_2_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3_1(253) WHEN s_2_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3_1(254) WHEN s_2_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3_1(255);

  
  out0_184 <= gmul2_1(0) WHEN s_1_1 = to_unsigned(16#01#, 8) ELSE
      gmul2_1(1) WHEN s_1_1 = to_unsigned(16#02#, 8) ELSE
      gmul2_1(2) WHEN s_1_1 = to_unsigned(16#03#, 8) ELSE
      gmul2_1(3) WHEN s_1_1 = to_unsigned(16#04#, 8) ELSE
      gmul2_1(4) WHEN s_1_1 = to_unsigned(16#05#, 8) ELSE
      gmul2_1(5) WHEN s_1_1 = to_unsigned(16#06#, 8) ELSE
      gmul2_1(6) WHEN s_1_1 = to_unsigned(16#07#, 8) ELSE
      gmul2_1(7) WHEN s_1_1 = to_unsigned(16#08#, 8) ELSE
      gmul2_1(8) WHEN s_1_1 = to_unsigned(16#09#, 8) ELSE
      gmul2_1(9) WHEN s_1_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2_1(10) WHEN s_1_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2_1(11) WHEN s_1_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2_1(12) WHEN s_1_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2_1(13) WHEN s_1_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2_1(14) WHEN s_1_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2_1(15) WHEN s_1_1 = to_unsigned(16#10#, 8) ELSE
      gmul2_1(16) WHEN s_1_1 = to_unsigned(16#11#, 8) ELSE
      gmul2_1(17) WHEN s_1_1 = to_unsigned(16#12#, 8) ELSE
      gmul2_1(18) WHEN s_1_1 = to_unsigned(16#13#, 8) ELSE
      gmul2_1(19) WHEN s_1_1 = to_unsigned(16#14#, 8) ELSE
      gmul2_1(20) WHEN s_1_1 = to_unsigned(16#15#, 8) ELSE
      gmul2_1(21) WHEN s_1_1 = to_unsigned(16#16#, 8) ELSE
      gmul2_1(22) WHEN s_1_1 = to_unsigned(16#17#, 8) ELSE
      gmul2_1(23) WHEN s_1_1 = to_unsigned(16#18#, 8) ELSE
      gmul2_1(24) WHEN s_1_1 = to_unsigned(16#19#, 8) ELSE
      gmul2_1(25) WHEN s_1_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2_1(26) WHEN s_1_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2_1(27) WHEN s_1_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2_1(28) WHEN s_1_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2_1(29) WHEN s_1_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2_1(30) WHEN s_1_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2_1(31) WHEN s_1_1 = to_unsigned(16#20#, 8) ELSE
      gmul2_1(32) WHEN s_1_1 = to_unsigned(16#21#, 8) ELSE
      gmul2_1(33) WHEN s_1_1 = to_unsigned(16#22#, 8) ELSE
      gmul2_1(34) WHEN s_1_1 = to_unsigned(16#23#, 8) ELSE
      gmul2_1(35) WHEN s_1_1 = to_unsigned(16#24#, 8) ELSE
      gmul2_1(36) WHEN s_1_1 = to_unsigned(16#25#, 8) ELSE
      gmul2_1(37) WHEN s_1_1 = to_unsigned(16#26#, 8) ELSE
      gmul2_1(38) WHEN s_1_1 = to_unsigned(16#27#, 8) ELSE
      gmul2_1(39) WHEN s_1_1 = to_unsigned(16#28#, 8) ELSE
      gmul2_1(40) WHEN s_1_1 = to_unsigned(16#29#, 8) ELSE
      gmul2_1(41) WHEN s_1_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2_1(42) WHEN s_1_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2_1(43) WHEN s_1_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2_1(44) WHEN s_1_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2_1(45) WHEN s_1_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2_1(46) WHEN s_1_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2_1(47) WHEN s_1_1 = to_unsigned(16#30#, 8) ELSE
      gmul2_1(48) WHEN s_1_1 = to_unsigned(16#31#, 8) ELSE
      gmul2_1(49) WHEN s_1_1 = to_unsigned(16#32#, 8) ELSE
      gmul2_1(50) WHEN s_1_1 = to_unsigned(16#33#, 8) ELSE
      gmul2_1(51) WHEN s_1_1 = to_unsigned(16#34#, 8) ELSE
      gmul2_1(52) WHEN s_1_1 = to_unsigned(16#35#, 8) ELSE
      gmul2_1(53) WHEN s_1_1 = to_unsigned(16#36#, 8) ELSE
      gmul2_1(54) WHEN s_1_1 = to_unsigned(16#37#, 8) ELSE
      gmul2_1(55) WHEN s_1_1 = to_unsigned(16#38#, 8) ELSE
      gmul2_1(56) WHEN s_1_1 = to_unsigned(16#39#, 8) ELSE
      gmul2_1(57) WHEN s_1_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2_1(58) WHEN s_1_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2_1(59) WHEN s_1_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2_1(60) WHEN s_1_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2_1(61) WHEN s_1_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2_1(62) WHEN s_1_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2_1(63) WHEN s_1_1 = to_unsigned(16#40#, 8) ELSE
      gmul2_1(64) WHEN s_1_1 = to_unsigned(16#41#, 8) ELSE
      gmul2_1(65) WHEN s_1_1 = to_unsigned(16#42#, 8) ELSE
      gmul2_1(66) WHEN s_1_1 = to_unsigned(16#43#, 8) ELSE
      gmul2_1(67) WHEN s_1_1 = to_unsigned(16#44#, 8) ELSE
      gmul2_1(68) WHEN s_1_1 = to_unsigned(16#45#, 8) ELSE
      gmul2_1(69) WHEN s_1_1 = to_unsigned(16#46#, 8) ELSE
      gmul2_1(70) WHEN s_1_1 = to_unsigned(16#47#, 8) ELSE
      gmul2_1(71) WHEN s_1_1 = to_unsigned(16#48#, 8) ELSE
      gmul2_1(72) WHEN s_1_1 = to_unsigned(16#49#, 8) ELSE
      gmul2_1(73) WHEN s_1_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2_1(74) WHEN s_1_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2_1(75) WHEN s_1_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2_1(76) WHEN s_1_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2_1(77) WHEN s_1_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2_1(78) WHEN s_1_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2_1(79) WHEN s_1_1 = to_unsigned(16#50#, 8) ELSE
      gmul2_1(80) WHEN s_1_1 = to_unsigned(16#51#, 8) ELSE
      gmul2_1(81) WHEN s_1_1 = to_unsigned(16#52#, 8) ELSE
      gmul2_1(82) WHEN s_1_1 = to_unsigned(16#53#, 8) ELSE
      gmul2_1(83) WHEN s_1_1 = to_unsigned(16#54#, 8) ELSE
      gmul2_1(84) WHEN s_1_1 = to_unsigned(16#55#, 8) ELSE
      gmul2_1(85) WHEN s_1_1 = to_unsigned(16#56#, 8) ELSE
      gmul2_1(86) WHEN s_1_1 = to_unsigned(16#57#, 8) ELSE
      gmul2_1(87) WHEN s_1_1 = to_unsigned(16#58#, 8) ELSE
      gmul2_1(88) WHEN s_1_1 = to_unsigned(16#59#, 8) ELSE
      gmul2_1(89) WHEN s_1_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2_1(90) WHEN s_1_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2_1(91) WHEN s_1_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2_1(92) WHEN s_1_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2_1(93) WHEN s_1_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2_1(94) WHEN s_1_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2_1(95) WHEN s_1_1 = to_unsigned(16#60#, 8) ELSE
      gmul2_1(96) WHEN s_1_1 = to_unsigned(16#61#, 8) ELSE
      gmul2_1(97) WHEN s_1_1 = to_unsigned(16#62#, 8) ELSE
      gmul2_1(98) WHEN s_1_1 = to_unsigned(16#63#, 8) ELSE
      gmul2_1(99) WHEN s_1_1 = to_unsigned(16#64#, 8) ELSE
      gmul2_1(100) WHEN s_1_1 = to_unsigned(16#65#, 8) ELSE
      gmul2_1(101) WHEN s_1_1 = to_unsigned(16#66#, 8) ELSE
      gmul2_1(102) WHEN s_1_1 = to_unsigned(16#67#, 8) ELSE
      gmul2_1(103) WHEN s_1_1 = to_unsigned(16#68#, 8) ELSE
      gmul2_1(104) WHEN s_1_1 = to_unsigned(16#69#, 8) ELSE
      gmul2_1(105) WHEN s_1_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2_1(106) WHEN s_1_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2_1(107) WHEN s_1_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2_1(108) WHEN s_1_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2_1(109) WHEN s_1_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2_1(110) WHEN s_1_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2_1(111) WHEN s_1_1 = to_unsigned(16#70#, 8) ELSE
      gmul2_1(112) WHEN s_1_1 = to_unsigned(16#71#, 8) ELSE
      gmul2_1(113) WHEN s_1_1 = to_unsigned(16#72#, 8) ELSE
      gmul2_1(114) WHEN s_1_1 = to_unsigned(16#73#, 8) ELSE
      gmul2_1(115) WHEN s_1_1 = to_unsigned(16#74#, 8) ELSE
      gmul2_1(116) WHEN s_1_1 = to_unsigned(16#75#, 8) ELSE
      gmul2_1(117) WHEN s_1_1 = to_unsigned(16#76#, 8) ELSE
      gmul2_1(118) WHEN s_1_1 = to_unsigned(16#77#, 8) ELSE
      gmul2_1(119) WHEN s_1_1 = to_unsigned(16#78#, 8) ELSE
      gmul2_1(120) WHEN s_1_1 = to_unsigned(16#79#, 8) ELSE
      gmul2_1(121) WHEN s_1_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2_1(122) WHEN s_1_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2_1(123) WHEN s_1_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2_1(124) WHEN s_1_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2_1(125) WHEN s_1_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2_1(126) WHEN s_1_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2_1(127) WHEN s_1_1 = to_unsigned(16#80#, 8) ELSE
      gmul2_1(128) WHEN s_1_1 = to_unsigned(16#81#, 8) ELSE
      gmul2_1(129) WHEN s_1_1 = to_unsigned(16#82#, 8) ELSE
      gmul2_1(130) WHEN s_1_1 = to_unsigned(16#83#, 8) ELSE
      gmul2_1(131) WHEN s_1_1 = to_unsigned(16#84#, 8) ELSE
      gmul2_1(132) WHEN s_1_1 = to_unsigned(16#85#, 8) ELSE
      gmul2_1(133) WHEN s_1_1 = to_unsigned(16#86#, 8) ELSE
      gmul2_1(134) WHEN s_1_1 = to_unsigned(16#87#, 8) ELSE
      gmul2_1(135) WHEN s_1_1 = to_unsigned(16#88#, 8) ELSE
      gmul2_1(136) WHEN s_1_1 = to_unsigned(16#89#, 8) ELSE
      gmul2_1(137) WHEN s_1_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2_1(138) WHEN s_1_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2_1(139) WHEN s_1_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2_1(140) WHEN s_1_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2_1(141) WHEN s_1_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2_1(142) WHEN s_1_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2_1(143) WHEN s_1_1 = to_unsigned(16#90#, 8) ELSE
      gmul2_1(144) WHEN s_1_1 = to_unsigned(16#91#, 8) ELSE
      gmul2_1(145) WHEN s_1_1 = to_unsigned(16#92#, 8) ELSE
      gmul2_1(146) WHEN s_1_1 = to_unsigned(16#93#, 8) ELSE
      gmul2_1(147) WHEN s_1_1 = to_unsigned(16#94#, 8) ELSE
      gmul2_1(148) WHEN s_1_1 = to_unsigned(16#95#, 8) ELSE
      gmul2_1(149) WHEN s_1_1 = to_unsigned(16#96#, 8) ELSE
      gmul2_1(150) WHEN s_1_1 = to_unsigned(16#97#, 8) ELSE
      gmul2_1(151) WHEN s_1_1 = to_unsigned(16#98#, 8) ELSE
      gmul2_1(152) WHEN s_1_1 = to_unsigned(16#99#, 8) ELSE
      gmul2_1(153) WHEN s_1_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2_1(154) WHEN s_1_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2_1(155) WHEN s_1_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2_1(156) WHEN s_1_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2_1(157) WHEN s_1_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2_1(158) WHEN s_1_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2_1(159) WHEN s_1_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2_1(160) WHEN s_1_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2_1(161) WHEN s_1_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2_1(162) WHEN s_1_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2_1(163) WHEN s_1_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2_1(164) WHEN s_1_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2_1(165) WHEN s_1_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2_1(166) WHEN s_1_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2_1(167) WHEN s_1_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2_1(168) WHEN s_1_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2_1(169) WHEN s_1_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2_1(170) WHEN s_1_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2_1(171) WHEN s_1_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2_1(172) WHEN s_1_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2_1(173) WHEN s_1_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2_1(174) WHEN s_1_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2_1(175) WHEN s_1_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2_1(176) WHEN s_1_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2_1(177) WHEN s_1_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2_1(178) WHEN s_1_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2_1(179) WHEN s_1_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2_1(180) WHEN s_1_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2_1(181) WHEN s_1_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2_1(182) WHEN s_1_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2_1(183) WHEN s_1_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2_1(184) WHEN s_1_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2_1(185) WHEN s_1_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2_1(186) WHEN s_1_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2_1(187) WHEN s_1_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2_1(188) WHEN s_1_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2_1(189) WHEN s_1_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2_1(190) WHEN s_1_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2_1(191) WHEN s_1_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2_1(192) WHEN s_1_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2_1(193) WHEN s_1_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2_1(194) WHEN s_1_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2_1(195) WHEN s_1_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2_1(196) WHEN s_1_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2_1(197) WHEN s_1_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2_1(198) WHEN s_1_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2_1(199) WHEN s_1_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2_1(200) WHEN s_1_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2_1(201) WHEN s_1_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2_1(202) WHEN s_1_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2_1(203) WHEN s_1_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2_1(204) WHEN s_1_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2_1(205) WHEN s_1_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2_1(206) WHEN s_1_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2_1(207) WHEN s_1_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2_1(208) WHEN s_1_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2_1(209) WHEN s_1_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2_1(210) WHEN s_1_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2_1(211) WHEN s_1_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2_1(212) WHEN s_1_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2_1(213) WHEN s_1_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2_1(214) WHEN s_1_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2_1(215) WHEN s_1_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2_1(216) WHEN s_1_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2_1(217) WHEN s_1_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2_1(218) WHEN s_1_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2_1(219) WHEN s_1_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2_1(220) WHEN s_1_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2_1(221) WHEN s_1_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2_1(222) WHEN s_1_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2_1(223) WHEN s_1_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2_1(224) WHEN s_1_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2_1(225) WHEN s_1_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2_1(226) WHEN s_1_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2_1(227) WHEN s_1_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2_1(228) WHEN s_1_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2_1(229) WHEN s_1_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2_1(230) WHEN s_1_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2_1(231) WHEN s_1_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2_1(232) WHEN s_1_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2_1(233) WHEN s_1_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2_1(234) WHEN s_1_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2_1(235) WHEN s_1_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2_1(236) WHEN s_1_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2_1(237) WHEN s_1_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2_1(238) WHEN s_1_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2_1(239) WHEN s_1_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2_1(240) WHEN s_1_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2_1(241) WHEN s_1_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2_1(242) WHEN s_1_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2_1(243) WHEN s_1_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2_1(244) WHEN s_1_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2_1(245) WHEN s_1_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2_1(246) WHEN s_1_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2_1(247) WHEN s_1_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2_1(248) WHEN s_1_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2_1(249) WHEN s_1_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2_1(250) WHEN s_1_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2_1(251) WHEN s_1_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2_1(252) WHEN s_1_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2_1(253) WHEN s_1_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2_1(254) WHEN s_1_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2_1(255);

  out0_185 <= s_0_1 XOR out0_184;

  b2_3 <= out0_185 XOR out0_183;

  out0_186 <= b2_3 XOR s_3_1;

  s_3_1 <= s_s_1(3);

  s_2_1 <= s_s_1(2);

  s_1_1 <= s_s_1(1);

  
  out0_187 <= gmul3(0) WHEN s_1_1 = to_unsigned(16#01#, 8) ELSE
      gmul3(1) WHEN s_1_1 = to_unsigned(16#02#, 8) ELSE
      gmul3(2) WHEN s_1_1 = to_unsigned(16#03#, 8) ELSE
      gmul3(3) WHEN s_1_1 = to_unsigned(16#04#, 8) ELSE
      gmul3(4) WHEN s_1_1 = to_unsigned(16#05#, 8) ELSE
      gmul3(5) WHEN s_1_1 = to_unsigned(16#06#, 8) ELSE
      gmul3(6) WHEN s_1_1 = to_unsigned(16#07#, 8) ELSE
      gmul3(7) WHEN s_1_1 = to_unsigned(16#08#, 8) ELSE
      gmul3(8) WHEN s_1_1 = to_unsigned(16#09#, 8) ELSE
      gmul3(9) WHEN s_1_1 = to_unsigned(16#0A#, 8) ELSE
      gmul3(10) WHEN s_1_1 = to_unsigned(16#0B#, 8) ELSE
      gmul3(11) WHEN s_1_1 = to_unsigned(16#0C#, 8) ELSE
      gmul3(12) WHEN s_1_1 = to_unsigned(16#0D#, 8) ELSE
      gmul3(13) WHEN s_1_1 = to_unsigned(16#0E#, 8) ELSE
      gmul3(14) WHEN s_1_1 = to_unsigned(16#0F#, 8) ELSE
      gmul3(15) WHEN s_1_1 = to_unsigned(16#10#, 8) ELSE
      gmul3(16) WHEN s_1_1 = to_unsigned(16#11#, 8) ELSE
      gmul3(17) WHEN s_1_1 = to_unsigned(16#12#, 8) ELSE
      gmul3(18) WHEN s_1_1 = to_unsigned(16#13#, 8) ELSE
      gmul3(19) WHEN s_1_1 = to_unsigned(16#14#, 8) ELSE
      gmul3(20) WHEN s_1_1 = to_unsigned(16#15#, 8) ELSE
      gmul3(21) WHEN s_1_1 = to_unsigned(16#16#, 8) ELSE
      gmul3(22) WHEN s_1_1 = to_unsigned(16#17#, 8) ELSE
      gmul3(23) WHEN s_1_1 = to_unsigned(16#18#, 8) ELSE
      gmul3(24) WHEN s_1_1 = to_unsigned(16#19#, 8) ELSE
      gmul3(25) WHEN s_1_1 = to_unsigned(16#1A#, 8) ELSE
      gmul3(26) WHEN s_1_1 = to_unsigned(16#1B#, 8) ELSE
      gmul3(27) WHEN s_1_1 = to_unsigned(16#1C#, 8) ELSE
      gmul3(28) WHEN s_1_1 = to_unsigned(16#1D#, 8) ELSE
      gmul3(29) WHEN s_1_1 = to_unsigned(16#1E#, 8) ELSE
      gmul3(30) WHEN s_1_1 = to_unsigned(16#1F#, 8) ELSE
      gmul3(31) WHEN s_1_1 = to_unsigned(16#20#, 8) ELSE
      gmul3(32) WHEN s_1_1 = to_unsigned(16#21#, 8) ELSE
      gmul3(33) WHEN s_1_1 = to_unsigned(16#22#, 8) ELSE
      gmul3(34) WHEN s_1_1 = to_unsigned(16#23#, 8) ELSE
      gmul3(35) WHEN s_1_1 = to_unsigned(16#24#, 8) ELSE
      gmul3(36) WHEN s_1_1 = to_unsigned(16#25#, 8) ELSE
      gmul3(37) WHEN s_1_1 = to_unsigned(16#26#, 8) ELSE
      gmul3(38) WHEN s_1_1 = to_unsigned(16#27#, 8) ELSE
      gmul3(39) WHEN s_1_1 = to_unsigned(16#28#, 8) ELSE
      gmul3(40) WHEN s_1_1 = to_unsigned(16#29#, 8) ELSE
      gmul3(41) WHEN s_1_1 = to_unsigned(16#2A#, 8) ELSE
      gmul3(42) WHEN s_1_1 = to_unsigned(16#2B#, 8) ELSE
      gmul3(43) WHEN s_1_1 = to_unsigned(16#2C#, 8) ELSE
      gmul3(44) WHEN s_1_1 = to_unsigned(16#2D#, 8) ELSE
      gmul3(45) WHEN s_1_1 = to_unsigned(16#2E#, 8) ELSE
      gmul3(46) WHEN s_1_1 = to_unsigned(16#2F#, 8) ELSE
      gmul3(47) WHEN s_1_1 = to_unsigned(16#30#, 8) ELSE
      gmul3(48) WHEN s_1_1 = to_unsigned(16#31#, 8) ELSE
      gmul3(49) WHEN s_1_1 = to_unsigned(16#32#, 8) ELSE
      gmul3(50) WHEN s_1_1 = to_unsigned(16#33#, 8) ELSE
      gmul3(51) WHEN s_1_1 = to_unsigned(16#34#, 8) ELSE
      gmul3(52) WHEN s_1_1 = to_unsigned(16#35#, 8) ELSE
      gmul3(53) WHEN s_1_1 = to_unsigned(16#36#, 8) ELSE
      gmul3(54) WHEN s_1_1 = to_unsigned(16#37#, 8) ELSE
      gmul3(55) WHEN s_1_1 = to_unsigned(16#38#, 8) ELSE
      gmul3(56) WHEN s_1_1 = to_unsigned(16#39#, 8) ELSE
      gmul3(57) WHEN s_1_1 = to_unsigned(16#3A#, 8) ELSE
      gmul3(58) WHEN s_1_1 = to_unsigned(16#3B#, 8) ELSE
      gmul3(59) WHEN s_1_1 = to_unsigned(16#3C#, 8) ELSE
      gmul3(60) WHEN s_1_1 = to_unsigned(16#3D#, 8) ELSE
      gmul3(61) WHEN s_1_1 = to_unsigned(16#3E#, 8) ELSE
      gmul3(62) WHEN s_1_1 = to_unsigned(16#3F#, 8) ELSE
      gmul3(63) WHEN s_1_1 = to_unsigned(16#40#, 8) ELSE
      gmul3(64) WHEN s_1_1 = to_unsigned(16#41#, 8) ELSE
      gmul3(65) WHEN s_1_1 = to_unsigned(16#42#, 8) ELSE
      gmul3(66) WHEN s_1_1 = to_unsigned(16#43#, 8) ELSE
      gmul3(67) WHEN s_1_1 = to_unsigned(16#44#, 8) ELSE
      gmul3(68) WHEN s_1_1 = to_unsigned(16#45#, 8) ELSE
      gmul3(69) WHEN s_1_1 = to_unsigned(16#46#, 8) ELSE
      gmul3(70) WHEN s_1_1 = to_unsigned(16#47#, 8) ELSE
      gmul3(71) WHEN s_1_1 = to_unsigned(16#48#, 8) ELSE
      gmul3(72) WHEN s_1_1 = to_unsigned(16#49#, 8) ELSE
      gmul3(73) WHEN s_1_1 = to_unsigned(16#4A#, 8) ELSE
      gmul3(74) WHEN s_1_1 = to_unsigned(16#4B#, 8) ELSE
      gmul3(75) WHEN s_1_1 = to_unsigned(16#4C#, 8) ELSE
      gmul3(76) WHEN s_1_1 = to_unsigned(16#4D#, 8) ELSE
      gmul3(77) WHEN s_1_1 = to_unsigned(16#4E#, 8) ELSE
      gmul3(78) WHEN s_1_1 = to_unsigned(16#4F#, 8) ELSE
      gmul3(79) WHEN s_1_1 = to_unsigned(16#50#, 8) ELSE
      gmul3(80) WHEN s_1_1 = to_unsigned(16#51#, 8) ELSE
      gmul3(81) WHEN s_1_1 = to_unsigned(16#52#, 8) ELSE
      gmul3(82) WHEN s_1_1 = to_unsigned(16#53#, 8) ELSE
      gmul3(83) WHEN s_1_1 = to_unsigned(16#54#, 8) ELSE
      gmul3(84) WHEN s_1_1 = to_unsigned(16#55#, 8) ELSE
      gmul3(85) WHEN s_1_1 = to_unsigned(16#56#, 8) ELSE
      gmul3(86) WHEN s_1_1 = to_unsigned(16#57#, 8) ELSE
      gmul3(87) WHEN s_1_1 = to_unsigned(16#58#, 8) ELSE
      gmul3(88) WHEN s_1_1 = to_unsigned(16#59#, 8) ELSE
      gmul3(89) WHEN s_1_1 = to_unsigned(16#5A#, 8) ELSE
      gmul3(90) WHEN s_1_1 = to_unsigned(16#5B#, 8) ELSE
      gmul3(91) WHEN s_1_1 = to_unsigned(16#5C#, 8) ELSE
      gmul3(92) WHEN s_1_1 = to_unsigned(16#5D#, 8) ELSE
      gmul3(93) WHEN s_1_1 = to_unsigned(16#5E#, 8) ELSE
      gmul3(94) WHEN s_1_1 = to_unsigned(16#5F#, 8) ELSE
      gmul3(95) WHEN s_1_1 = to_unsigned(16#60#, 8) ELSE
      gmul3(96) WHEN s_1_1 = to_unsigned(16#61#, 8) ELSE
      gmul3(97) WHEN s_1_1 = to_unsigned(16#62#, 8) ELSE
      gmul3(98) WHEN s_1_1 = to_unsigned(16#63#, 8) ELSE
      gmul3(99) WHEN s_1_1 = to_unsigned(16#64#, 8) ELSE
      gmul3(100) WHEN s_1_1 = to_unsigned(16#65#, 8) ELSE
      gmul3(101) WHEN s_1_1 = to_unsigned(16#66#, 8) ELSE
      gmul3(102) WHEN s_1_1 = to_unsigned(16#67#, 8) ELSE
      gmul3(103) WHEN s_1_1 = to_unsigned(16#68#, 8) ELSE
      gmul3(104) WHEN s_1_1 = to_unsigned(16#69#, 8) ELSE
      gmul3(105) WHEN s_1_1 = to_unsigned(16#6A#, 8) ELSE
      gmul3(106) WHEN s_1_1 = to_unsigned(16#6B#, 8) ELSE
      gmul3(107) WHEN s_1_1 = to_unsigned(16#6C#, 8) ELSE
      gmul3(108) WHEN s_1_1 = to_unsigned(16#6D#, 8) ELSE
      gmul3(109) WHEN s_1_1 = to_unsigned(16#6E#, 8) ELSE
      gmul3(110) WHEN s_1_1 = to_unsigned(16#6F#, 8) ELSE
      gmul3(111) WHEN s_1_1 = to_unsigned(16#70#, 8) ELSE
      gmul3(112) WHEN s_1_1 = to_unsigned(16#71#, 8) ELSE
      gmul3(113) WHEN s_1_1 = to_unsigned(16#72#, 8) ELSE
      gmul3(114) WHEN s_1_1 = to_unsigned(16#73#, 8) ELSE
      gmul3(115) WHEN s_1_1 = to_unsigned(16#74#, 8) ELSE
      gmul3(116) WHEN s_1_1 = to_unsigned(16#75#, 8) ELSE
      gmul3(117) WHEN s_1_1 = to_unsigned(16#76#, 8) ELSE
      gmul3(118) WHEN s_1_1 = to_unsigned(16#77#, 8) ELSE
      gmul3(119) WHEN s_1_1 = to_unsigned(16#78#, 8) ELSE
      gmul3(120) WHEN s_1_1 = to_unsigned(16#79#, 8) ELSE
      gmul3(121) WHEN s_1_1 = to_unsigned(16#7A#, 8) ELSE
      gmul3(122) WHEN s_1_1 = to_unsigned(16#7B#, 8) ELSE
      gmul3(123) WHEN s_1_1 = to_unsigned(16#7C#, 8) ELSE
      gmul3(124) WHEN s_1_1 = to_unsigned(16#7D#, 8) ELSE
      gmul3(125) WHEN s_1_1 = to_unsigned(16#7E#, 8) ELSE
      gmul3(126) WHEN s_1_1 = to_unsigned(16#7F#, 8) ELSE
      gmul3(127) WHEN s_1_1 = to_unsigned(16#80#, 8) ELSE
      gmul3(128) WHEN s_1_1 = to_unsigned(16#81#, 8) ELSE
      gmul3(129) WHEN s_1_1 = to_unsigned(16#82#, 8) ELSE
      gmul3(130) WHEN s_1_1 = to_unsigned(16#83#, 8) ELSE
      gmul3(131) WHEN s_1_1 = to_unsigned(16#84#, 8) ELSE
      gmul3(132) WHEN s_1_1 = to_unsigned(16#85#, 8) ELSE
      gmul3(133) WHEN s_1_1 = to_unsigned(16#86#, 8) ELSE
      gmul3(134) WHEN s_1_1 = to_unsigned(16#87#, 8) ELSE
      gmul3(135) WHEN s_1_1 = to_unsigned(16#88#, 8) ELSE
      gmul3(136) WHEN s_1_1 = to_unsigned(16#89#, 8) ELSE
      gmul3(137) WHEN s_1_1 = to_unsigned(16#8A#, 8) ELSE
      gmul3(138) WHEN s_1_1 = to_unsigned(16#8B#, 8) ELSE
      gmul3(139) WHEN s_1_1 = to_unsigned(16#8C#, 8) ELSE
      gmul3(140) WHEN s_1_1 = to_unsigned(16#8D#, 8) ELSE
      gmul3(141) WHEN s_1_1 = to_unsigned(16#8E#, 8) ELSE
      gmul3(142) WHEN s_1_1 = to_unsigned(16#8F#, 8) ELSE
      gmul3(143) WHEN s_1_1 = to_unsigned(16#90#, 8) ELSE
      gmul3(144) WHEN s_1_1 = to_unsigned(16#91#, 8) ELSE
      gmul3(145) WHEN s_1_1 = to_unsigned(16#92#, 8) ELSE
      gmul3(146) WHEN s_1_1 = to_unsigned(16#93#, 8) ELSE
      gmul3(147) WHEN s_1_1 = to_unsigned(16#94#, 8) ELSE
      gmul3(148) WHEN s_1_1 = to_unsigned(16#95#, 8) ELSE
      gmul3(149) WHEN s_1_1 = to_unsigned(16#96#, 8) ELSE
      gmul3(150) WHEN s_1_1 = to_unsigned(16#97#, 8) ELSE
      gmul3(151) WHEN s_1_1 = to_unsigned(16#98#, 8) ELSE
      gmul3(152) WHEN s_1_1 = to_unsigned(16#99#, 8) ELSE
      gmul3(153) WHEN s_1_1 = to_unsigned(16#9A#, 8) ELSE
      gmul3(154) WHEN s_1_1 = to_unsigned(16#9B#, 8) ELSE
      gmul3(155) WHEN s_1_1 = to_unsigned(16#9C#, 8) ELSE
      gmul3(156) WHEN s_1_1 = to_unsigned(16#9D#, 8) ELSE
      gmul3(157) WHEN s_1_1 = to_unsigned(16#9E#, 8) ELSE
      gmul3(158) WHEN s_1_1 = to_unsigned(16#9F#, 8) ELSE
      gmul3(159) WHEN s_1_1 = to_unsigned(16#A0#, 8) ELSE
      gmul3(160) WHEN s_1_1 = to_unsigned(16#A1#, 8) ELSE
      gmul3(161) WHEN s_1_1 = to_unsigned(16#A2#, 8) ELSE
      gmul3(162) WHEN s_1_1 = to_unsigned(16#A3#, 8) ELSE
      gmul3(163) WHEN s_1_1 = to_unsigned(16#A4#, 8) ELSE
      gmul3(164) WHEN s_1_1 = to_unsigned(16#A5#, 8) ELSE
      gmul3(165) WHEN s_1_1 = to_unsigned(16#A6#, 8) ELSE
      gmul3(166) WHEN s_1_1 = to_unsigned(16#A7#, 8) ELSE
      gmul3(167) WHEN s_1_1 = to_unsigned(16#A8#, 8) ELSE
      gmul3(168) WHEN s_1_1 = to_unsigned(16#A9#, 8) ELSE
      gmul3(169) WHEN s_1_1 = to_unsigned(16#AA#, 8) ELSE
      gmul3(170) WHEN s_1_1 = to_unsigned(16#AB#, 8) ELSE
      gmul3(171) WHEN s_1_1 = to_unsigned(16#AC#, 8) ELSE
      gmul3(172) WHEN s_1_1 = to_unsigned(16#AD#, 8) ELSE
      gmul3(173) WHEN s_1_1 = to_unsigned(16#AE#, 8) ELSE
      gmul3(174) WHEN s_1_1 = to_unsigned(16#AF#, 8) ELSE
      gmul3(175) WHEN s_1_1 = to_unsigned(16#B0#, 8) ELSE
      gmul3(176) WHEN s_1_1 = to_unsigned(16#B1#, 8) ELSE
      gmul3(177) WHEN s_1_1 = to_unsigned(16#B2#, 8) ELSE
      gmul3(178) WHEN s_1_1 = to_unsigned(16#B3#, 8) ELSE
      gmul3(179) WHEN s_1_1 = to_unsigned(16#B4#, 8) ELSE
      gmul3(180) WHEN s_1_1 = to_unsigned(16#B5#, 8) ELSE
      gmul3(181) WHEN s_1_1 = to_unsigned(16#B6#, 8) ELSE
      gmul3(182) WHEN s_1_1 = to_unsigned(16#B7#, 8) ELSE
      gmul3(183) WHEN s_1_1 = to_unsigned(16#B8#, 8) ELSE
      gmul3(184) WHEN s_1_1 = to_unsigned(16#B9#, 8) ELSE
      gmul3(185) WHEN s_1_1 = to_unsigned(16#BA#, 8) ELSE
      gmul3(186) WHEN s_1_1 = to_unsigned(16#BB#, 8) ELSE
      gmul3(187) WHEN s_1_1 = to_unsigned(16#BC#, 8) ELSE
      gmul3(188) WHEN s_1_1 = to_unsigned(16#BD#, 8) ELSE
      gmul3(189) WHEN s_1_1 = to_unsigned(16#BE#, 8) ELSE
      gmul3(190) WHEN s_1_1 = to_unsigned(16#BF#, 8) ELSE
      gmul3(191) WHEN s_1_1 = to_unsigned(16#C0#, 8) ELSE
      gmul3(192) WHEN s_1_1 = to_unsigned(16#C1#, 8) ELSE
      gmul3(193) WHEN s_1_1 = to_unsigned(16#C2#, 8) ELSE
      gmul3(194) WHEN s_1_1 = to_unsigned(16#C3#, 8) ELSE
      gmul3(195) WHEN s_1_1 = to_unsigned(16#C4#, 8) ELSE
      gmul3(196) WHEN s_1_1 = to_unsigned(16#C5#, 8) ELSE
      gmul3(197) WHEN s_1_1 = to_unsigned(16#C6#, 8) ELSE
      gmul3(198) WHEN s_1_1 = to_unsigned(16#C7#, 8) ELSE
      gmul3(199) WHEN s_1_1 = to_unsigned(16#C8#, 8) ELSE
      gmul3(200) WHEN s_1_1 = to_unsigned(16#C9#, 8) ELSE
      gmul3(201) WHEN s_1_1 = to_unsigned(16#CA#, 8) ELSE
      gmul3(202) WHEN s_1_1 = to_unsigned(16#CB#, 8) ELSE
      gmul3(203) WHEN s_1_1 = to_unsigned(16#CC#, 8) ELSE
      gmul3(204) WHEN s_1_1 = to_unsigned(16#CD#, 8) ELSE
      gmul3(205) WHEN s_1_1 = to_unsigned(16#CE#, 8) ELSE
      gmul3(206) WHEN s_1_1 = to_unsigned(16#CF#, 8) ELSE
      gmul3(207) WHEN s_1_1 = to_unsigned(16#D0#, 8) ELSE
      gmul3(208) WHEN s_1_1 = to_unsigned(16#D1#, 8) ELSE
      gmul3(209) WHEN s_1_1 = to_unsigned(16#D2#, 8) ELSE
      gmul3(210) WHEN s_1_1 = to_unsigned(16#D3#, 8) ELSE
      gmul3(211) WHEN s_1_1 = to_unsigned(16#D4#, 8) ELSE
      gmul3(212) WHEN s_1_1 = to_unsigned(16#D5#, 8) ELSE
      gmul3(213) WHEN s_1_1 = to_unsigned(16#D6#, 8) ELSE
      gmul3(214) WHEN s_1_1 = to_unsigned(16#D7#, 8) ELSE
      gmul3(215) WHEN s_1_1 = to_unsigned(16#D8#, 8) ELSE
      gmul3(216) WHEN s_1_1 = to_unsigned(16#D9#, 8) ELSE
      gmul3(217) WHEN s_1_1 = to_unsigned(16#DA#, 8) ELSE
      gmul3(218) WHEN s_1_1 = to_unsigned(16#DB#, 8) ELSE
      gmul3(219) WHEN s_1_1 = to_unsigned(16#DC#, 8) ELSE
      gmul3(220) WHEN s_1_1 = to_unsigned(16#DD#, 8) ELSE
      gmul3(221) WHEN s_1_1 = to_unsigned(16#DE#, 8) ELSE
      gmul3(222) WHEN s_1_1 = to_unsigned(16#DF#, 8) ELSE
      gmul3(223) WHEN s_1_1 = to_unsigned(16#E0#, 8) ELSE
      gmul3(224) WHEN s_1_1 = to_unsigned(16#E1#, 8) ELSE
      gmul3(225) WHEN s_1_1 = to_unsigned(16#E2#, 8) ELSE
      gmul3(226) WHEN s_1_1 = to_unsigned(16#E3#, 8) ELSE
      gmul3(227) WHEN s_1_1 = to_unsigned(16#E4#, 8) ELSE
      gmul3(228) WHEN s_1_1 = to_unsigned(16#E5#, 8) ELSE
      gmul3(229) WHEN s_1_1 = to_unsigned(16#E6#, 8) ELSE
      gmul3(230) WHEN s_1_1 = to_unsigned(16#E7#, 8) ELSE
      gmul3(231) WHEN s_1_1 = to_unsigned(16#E8#, 8) ELSE
      gmul3(232) WHEN s_1_1 = to_unsigned(16#E9#, 8) ELSE
      gmul3(233) WHEN s_1_1 = to_unsigned(16#EA#, 8) ELSE
      gmul3(234) WHEN s_1_1 = to_unsigned(16#EB#, 8) ELSE
      gmul3(235) WHEN s_1_1 = to_unsigned(16#EC#, 8) ELSE
      gmul3(236) WHEN s_1_1 = to_unsigned(16#ED#, 8) ELSE
      gmul3(237) WHEN s_1_1 = to_unsigned(16#EE#, 8) ELSE
      gmul3(238) WHEN s_1_1 = to_unsigned(16#EF#, 8) ELSE
      gmul3(239) WHEN s_1_1 = to_unsigned(16#F0#, 8) ELSE
      gmul3(240) WHEN s_1_1 = to_unsigned(16#F1#, 8) ELSE
      gmul3(241) WHEN s_1_1 = to_unsigned(16#F2#, 8) ELSE
      gmul3(242) WHEN s_1_1 = to_unsigned(16#F3#, 8) ELSE
      gmul3(243) WHEN s_1_1 = to_unsigned(16#F4#, 8) ELSE
      gmul3(244) WHEN s_1_1 = to_unsigned(16#F5#, 8) ELSE
      gmul3(245) WHEN s_1_1 = to_unsigned(16#F6#, 8) ELSE
      gmul3(246) WHEN s_1_1 = to_unsigned(16#F7#, 8) ELSE
      gmul3(247) WHEN s_1_1 = to_unsigned(16#F8#, 8) ELSE
      gmul3(248) WHEN s_1_1 = to_unsigned(16#F9#, 8) ELSE
      gmul3(249) WHEN s_1_1 = to_unsigned(16#FA#, 8) ELSE
      gmul3(250) WHEN s_1_1 = to_unsigned(16#FB#, 8) ELSE
      gmul3(251) WHEN s_1_1 = to_unsigned(16#FC#, 8) ELSE
      gmul3(252) WHEN s_1_1 = to_unsigned(16#FD#, 8) ELSE
      gmul3(253) WHEN s_1_1 = to_unsigned(16#FE#, 8) ELSE
      gmul3(254) WHEN s_1_1 = to_unsigned(16#FF#, 8) ELSE
      gmul3(255);

  s_0_1 <= s_s_1(0);

  
  out0_188 <= gmul2(0) WHEN s_0_1 = to_unsigned(16#01#, 8) ELSE
      gmul2(1) WHEN s_0_1 = to_unsigned(16#02#, 8) ELSE
      gmul2(2) WHEN s_0_1 = to_unsigned(16#03#, 8) ELSE
      gmul2(3) WHEN s_0_1 = to_unsigned(16#04#, 8) ELSE
      gmul2(4) WHEN s_0_1 = to_unsigned(16#05#, 8) ELSE
      gmul2(5) WHEN s_0_1 = to_unsigned(16#06#, 8) ELSE
      gmul2(6) WHEN s_0_1 = to_unsigned(16#07#, 8) ELSE
      gmul2(7) WHEN s_0_1 = to_unsigned(16#08#, 8) ELSE
      gmul2(8) WHEN s_0_1 = to_unsigned(16#09#, 8) ELSE
      gmul2(9) WHEN s_0_1 = to_unsigned(16#0A#, 8) ELSE
      gmul2(10) WHEN s_0_1 = to_unsigned(16#0B#, 8) ELSE
      gmul2(11) WHEN s_0_1 = to_unsigned(16#0C#, 8) ELSE
      gmul2(12) WHEN s_0_1 = to_unsigned(16#0D#, 8) ELSE
      gmul2(13) WHEN s_0_1 = to_unsigned(16#0E#, 8) ELSE
      gmul2(14) WHEN s_0_1 = to_unsigned(16#0F#, 8) ELSE
      gmul2(15) WHEN s_0_1 = to_unsigned(16#10#, 8) ELSE
      gmul2(16) WHEN s_0_1 = to_unsigned(16#11#, 8) ELSE
      gmul2(17) WHEN s_0_1 = to_unsigned(16#12#, 8) ELSE
      gmul2(18) WHEN s_0_1 = to_unsigned(16#13#, 8) ELSE
      gmul2(19) WHEN s_0_1 = to_unsigned(16#14#, 8) ELSE
      gmul2(20) WHEN s_0_1 = to_unsigned(16#15#, 8) ELSE
      gmul2(21) WHEN s_0_1 = to_unsigned(16#16#, 8) ELSE
      gmul2(22) WHEN s_0_1 = to_unsigned(16#17#, 8) ELSE
      gmul2(23) WHEN s_0_1 = to_unsigned(16#18#, 8) ELSE
      gmul2(24) WHEN s_0_1 = to_unsigned(16#19#, 8) ELSE
      gmul2(25) WHEN s_0_1 = to_unsigned(16#1A#, 8) ELSE
      gmul2(26) WHEN s_0_1 = to_unsigned(16#1B#, 8) ELSE
      gmul2(27) WHEN s_0_1 = to_unsigned(16#1C#, 8) ELSE
      gmul2(28) WHEN s_0_1 = to_unsigned(16#1D#, 8) ELSE
      gmul2(29) WHEN s_0_1 = to_unsigned(16#1E#, 8) ELSE
      gmul2(30) WHEN s_0_1 = to_unsigned(16#1F#, 8) ELSE
      gmul2(31) WHEN s_0_1 = to_unsigned(16#20#, 8) ELSE
      gmul2(32) WHEN s_0_1 = to_unsigned(16#21#, 8) ELSE
      gmul2(33) WHEN s_0_1 = to_unsigned(16#22#, 8) ELSE
      gmul2(34) WHEN s_0_1 = to_unsigned(16#23#, 8) ELSE
      gmul2(35) WHEN s_0_1 = to_unsigned(16#24#, 8) ELSE
      gmul2(36) WHEN s_0_1 = to_unsigned(16#25#, 8) ELSE
      gmul2(37) WHEN s_0_1 = to_unsigned(16#26#, 8) ELSE
      gmul2(38) WHEN s_0_1 = to_unsigned(16#27#, 8) ELSE
      gmul2(39) WHEN s_0_1 = to_unsigned(16#28#, 8) ELSE
      gmul2(40) WHEN s_0_1 = to_unsigned(16#29#, 8) ELSE
      gmul2(41) WHEN s_0_1 = to_unsigned(16#2A#, 8) ELSE
      gmul2(42) WHEN s_0_1 = to_unsigned(16#2B#, 8) ELSE
      gmul2(43) WHEN s_0_1 = to_unsigned(16#2C#, 8) ELSE
      gmul2(44) WHEN s_0_1 = to_unsigned(16#2D#, 8) ELSE
      gmul2(45) WHEN s_0_1 = to_unsigned(16#2E#, 8) ELSE
      gmul2(46) WHEN s_0_1 = to_unsigned(16#2F#, 8) ELSE
      gmul2(47) WHEN s_0_1 = to_unsigned(16#30#, 8) ELSE
      gmul2(48) WHEN s_0_1 = to_unsigned(16#31#, 8) ELSE
      gmul2(49) WHEN s_0_1 = to_unsigned(16#32#, 8) ELSE
      gmul2(50) WHEN s_0_1 = to_unsigned(16#33#, 8) ELSE
      gmul2(51) WHEN s_0_1 = to_unsigned(16#34#, 8) ELSE
      gmul2(52) WHEN s_0_1 = to_unsigned(16#35#, 8) ELSE
      gmul2(53) WHEN s_0_1 = to_unsigned(16#36#, 8) ELSE
      gmul2(54) WHEN s_0_1 = to_unsigned(16#37#, 8) ELSE
      gmul2(55) WHEN s_0_1 = to_unsigned(16#38#, 8) ELSE
      gmul2(56) WHEN s_0_1 = to_unsigned(16#39#, 8) ELSE
      gmul2(57) WHEN s_0_1 = to_unsigned(16#3A#, 8) ELSE
      gmul2(58) WHEN s_0_1 = to_unsigned(16#3B#, 8) ELSE
      gmul2(59) WHEN s_0_1 = to_unsigned(16#3C#, 8) ELSE
      gmul2(60) WHEN s_0_1 = to_unsigned(16#3D#, 8) ELSE
      gmul2(61) WHEN s_0_1 = to_unsigned(16#3E#, 8) ELSE
      gmul2(62) WHEN s_0_1 = to_unsigned(16#3F#, 8) ELSE
      gmul2(63) WHEN s_0_1 = to_unsigned(16#40#, 8) ELSE
      gmul2(64) WHEN s_0_1 = to_unsigned(16#41#, 8) ELSE
      gmul2(65) WHEN s_0_1 = to_unsigned(16#42#, 8) ELSE
      gmul2(66) WHEN s_0_1 = to_unsigned(16#43#, 8) ELSE
      gmul2(67) WHEN s_0_1 = to_unsigned(16#44#, 8) ELSE
      gmul2(68) WHEN s_0_1 = to_unsigned(16#45#, 8) ELSE
      gmul2(69) WHEN s_0_1 = to_unsigned(16#46#, 8) ELSE
      gmul2(70) WHEN s_0_1 = to_unsigned(16#47#, 8) ELSE
      gmul2(71) WHEN s_0_1 = to_unsigned(16#48#, 8) ELSE
      gmul2(72) WHEN s_0_1 = to_unsigned(16#49#, 8) ELSE
      gmul2(73) WHEN s_0_1 = to_unsigned(16#4A#, 8) ELSE
      gmul2(74) WHEN s_0_1 = to_unsigned(16#4B#, 8) ELSE
      gmul2(75) WHEN s_0_1 = to_unsigned(16#4C#, 8) ELSE
      gmul2(76) WHEN s_0_1 = to_unsigned(16#4D#, 8) ELSE
      gmul2(77) WHEN s_0_1 = to_unsigned(16#4E#, 8) ELSE
      gmul2(78) WHEN s_0_1 = to_unsigned(16#4F#, 8) ELSE
      gmul2(79) WHEN s_0_1 = to_unsigned(16#50#, 8) ELSE
      gmul2(80) WHEN s_0_1 = to_unsigned(16#51#, 8) ELSE
      gmul2(81) WHEN s_0_1 = to_unsigned(16#52#, 8) ELSE
      gmul2(82) WHEN s_0_1 = to_unsigned(16#53#, 8) ELSE
      gmul2(83) WHEN s_0_1 = to_unsigned(16#54#, 8) ELSE
      gmul2(84) WHEN s_0_1 = to_unsigned(16#55#, 8) ELSE
      gmul2(85) WHEN s_0_1 = to_unsigned(16#56#, 8) ELSE
      gmul2(86) WHEN s_0_1 = to_unsigned(16#57#, 8) ELSE
      gmul2(87) WHEN s_0_1 = to_unsigned(16#58#, 8) ELSE
      gmul2(88) WHEN s_0_1 = to_unsigned(16#59#, 8) ELSE
      gmul2(89) WHEN s_0_1 = to_unsigned(16#5A#, 8) ELSE
      gmul2(90) WHEN s_0_1 = to_unsigned(16#5B#, 8) ELSE
      gmul2(91) WHEN s_0_1 = to_unsigned(16#5C#, 8) ELSE
      gmul2(92) WHEN s_0_1 = to_unsigned(16#5D#, 8) ELSE
      gmul2(93) WHEN s_0_1 = to_unsigned(16#5E#, 8) ELSE
      gmul2(94) WHEN s_0_1 = to_unsigned(16#5F#, 8) ELSE
      gmul2(95) WHEN s_0_1 = to_unsigned(16#60#, 8) ELSE
      gmul2(96) WHEN s_0_1 = to_unsigned(16#61#, 8) ELSE
      gmul2(97) WHEN s_0_1 = to_unsigned(16#62#, 8) ELSE
      gmul2(98) WHEN s_0_1 = to_unsigned(16#63#, 8) ELSE
      gmul2(99) WHEN s_0_1 = to_unsigned(16#64#, 8) ELSE
      gmul2(100) WHEN s_0_1 = to_unsigned(16#65#, 8) ELSE
      gmul2(101) WHEN s_0_1 = to_unsigned(16#66#, 8) ELSE
      gmul2(102) WHEN s_0_1 = to_unsigned(16#67#, 8) ELSE
      gmul2(103) WHEN s_0_1 = to_unsigned(16#68#, 8) ELSE
      gmul2(104) WHEN s_0_1 = to_unsigned(16#69#, 8) ELSE
      gmul2(105) WHEN s_0_1 = to_unsigned(16#6A#, 8) ELSE
      gmul2(106) WHEN s_0_1 = to_unsigned(16#6B#, 8) ELSE
      gmul2(107) WHEN s_0_1 = to_unsigned(16#6C#, 8) ELSE
      gmul2(108) WHEN s_0_1 = to_unsigned(16#6D#, 8) ELSE
      gmul2(109) WHEN s_0_1 = to_unsigned(16#6E#, 8) ELSE
      gmul2(110) WHEN s_0_1 = to_unsigned(16#6F#, 8) ELSE
      gmul2(111) WHEN s_0_1 = to_unsigned(16#70#, 8) ELSE
      gmul2(112) WHEN s_0_1 = to_unsigned(16#71#, 8) ELSE
      gmul2(113) WHEN s_0_1 = to_unsigned(16#72#, 8) ELSE
      gmul2(114) WHEN s_0_1 = to_unsigned(16#73#, 8) ELSE
      gmul2(115) WHEN s_0_1 = to_unsigned(16#74#, 8) ELSE
      gmul2(116) WHEN s_0_1 = to_unsigned(16#75#, 8) ELSE
      gmul2(117) WHEN s_0_1 = to_unsigned(16#76#, 8) ELSE
      gmul2(118) WHEN s_0_1 = to_unsigned(16#77#, 8) ELSE
      gmul2(119) WHEN s_0_1 = to_unsigned(16#78#, 8) ELSE
      gmul2(120) WHEN s_0_1 = to_unsigned(16#79#, 8) ELSE
      gmul2(121) WHEN s_0_1 = to_unsigned(16#7A#, 8) ELSE
      gmul2(122) WHEN s_0_1 = to_unsigned(16#7B#, 8) ELSE
      gmul2(123) WHEN s_0_1 = to_unsigned(16#7C#, 8) ELSE
      gmul2(124) WHEN s_0_1 = to_unsigned(16#7D#, 8) ELSE
      gmul2(125) WHEN s_0_1 = to_unsigned(16#7E#, 8) ELSE
      gmul2(126) WHEN s_0_1 = to_unsigned(16#7F#, 8) ELSE
      gmul2(127) WHEN s_0_1 = to_unsigned(16#80#, 8) ELSE
      gmul2(128) WHEN s_0_1 = to_unsigned(16#81#, 8) ELSE
      gmul2(129) WHEN s_0_1 = to_unsigned(16#82#, 8) ELSE
      gmul2(130) WHEN s_0_1 = to_unsigned(16#83#, 8) ELSE
      gmul2(131) WHEN s_0_1 = to_unsigned(16#84#, 8) ELSE
      gmul2(132) WHEN s_0_1 = to_unsigned(16#85#, 8) ELSE
      gmul2(133) WHEN s_0_1 = to_unsigned(16#86#, 8) ELSE
      gmul2(134) WHEN s_0_1 = to_unsigned(16#87#, 8) ELSE
      gmul2(135) WHEN s_0_1 = to_unsigned(16#88#, 8) ELSE
      gmul2(136) WHEN s_0_1 = to_unsigned(16#89#, 8) ELSE
      gmul2(137) WHEN s_0_1 = to_unsigned(16#8A#, 8) ELSE
      gmul2(138) WHEN s_0_1 = to_unsigned(16#8B#, 8) ELSE
      gmul2(139) WHEN s_0_1 = to_unsigned(16#8C#, 8) ELSE
      gmul2(140) WHEN s_0_1 = to_unsigned(16#8D#, 8) ELSE
      gmul2(141) WHEN s_0_1 = to_unsigned(16#8E#, 8) ELSE
      gmul2(142) WHEN s_0_1 = to_unsigned(16#8F#, 8) ELSE
      gmul2(143) WHEN s_0_1 = to_unsigned(16#90#, 8) ELSE
      gmul2(144) WHEN s_0_1 = to_unsigned(16#91#, 8) ELSE
      gmul2(145) WHEN s_0_1 = to_unsigned(16#92#, 8) ELSE
      gmul2(146) WHEN s_0_1 = to_unsigned(16#93#, 8) ELSE
      gmul2(147) WHEN s_0_1 = to_unsigned(16#94#, 8) ELSE
      gmul2(148) WHEN s_0_1 = to_unsigned(16#95#, 8) ELSE
      gmul2(149) WHEN s_0_1 = to_unsigned(16#96#, 8) ELSE
      gmul2(150) WHEN s_0_1 = to_unsigned(16#97#, 8) ELSE
      gmul2(151) WHEN s_0_1 = to_unsigned(16#98#, 8) ELSE
      gmul2(152) WHEN s_0_1 = to_unsigned(16#99#, 8) ELSE
      gmul2(153) WHEN s_0_1 = to_unsigned(16#9A#, 8) ELSE
      gmul2(154) WHEN s_0_1 = to_unsigned(16#9B#, 8) ELSE
      gmul2(155) WHEN s_0_1 = to_unsigned(16#9C#, 8) ELSE
      gmul2(156) WHEN s_0_1 = to_unsigned(16#9D#, 8) ELSE
      gmul2(157) WHEN s_0_1 = to_unsigned(16#9E#, 8) ELSE
      gmul2(158) WHEN s_0_1 = to_unsigned(16#9F#, 8) ELSE
      gmul2(159) WHEN s_0_1 = to_unsigned(16#A0#, 8) ELSE
      gmul2(160) WHEN s_0_1 = to_unsigned(16#A1#, 8) ELSE
      gmul2(161) WHEN s_0_1 = to_unsigned(16#A2#, 8) ELSE
      gmul2(162) WHEN s_0_1 = to_unsigned(16#A3#, 8) ELSE
      gmul2(163) WHEN s_0_1 = to_unsigned(16#A4#, 8) ELSE
      gmul2(164) WHEN s_0_1 = to_unsigned(16#A5#, 8) ELSE
      gmul2(165) WHEN s_0_1 = to_unsigned(16#A6#, 8) ELSE
      gmul2(166) WHEN s_0_1 = to_unsigned(16#A7#, 8) ELSE
      gmul2(167) WHEN s_0_1 = to_unsigned(16#A8#, 8) ELSE
      gmul2(168) WHEN s_0_1 = to_unsigned(16#A9#, 8) ELSE
      gmul2(169) WHEN s_0_1 = to_unsigned(16#AA#, 8) ELSE
      gmul2(170) WHEN s_0_1 = to_unsigned(16#AB#, 8) ELSE
      gmul2(171) WHEN s_0_1 = to_unsigned(16#AC#, 8) ELSE
      gmul2(172) WHEN s_0_1 = to_unsigned(16#AD#, 8) ELSE
      gmul2(173) WHEN s_0_1 = to_unsigned(16#AE#, 8) ELSE
      gmul2(174) WHEN s_0_1 = to_unsigned(16#AF#, 8) ELSE
      gmul2(175) WHEN s_0_1 = to_unsigned(16#B0#, 8) ELSE
      gmul2(176) WHEN s_0_1 = to_unsigned(16#B1#, 8) ELSE
      gmul2(177) WHEN s_0_1 = to_unsigned(16#B2#, 8) ELSE
      gmul2(178) WHEN s_0_1 = to_unsigned(16#B3#, 8) ELSE
      gmul2(179) WHEN s_0_1 = to_unsigned(16#B4#, 8) ELSE
      gmul2(180) WHEN s_0_1 = to_unsigned(16#B5#, 8) ELSE
      gmul2(181) WHEN s_0_1 = to_unsigned(16#B6#, 8) ELSE
      gmul2(182) WHEN s_0_1 = to_unsigned(16#B7#, 8) ELSE
      gmul2(183) WHEN s_0_1 = to_unsigned(16#B8#, 8) ELSE
      gmul2(184) WHEN s_0_1 = to_unsigned(16#B9#, 8) ELSE
      gmul2(185) WHEN s_0_1 = to_unsigned(16#BA#, 8) ELSE
      gmul2(186) WHEN s_0_1 = to_unsigned(16#BB#, 8) ELSE
      gmul2(187) WHEN s_0_1 = to_unsigned(16#BC#, 8) ELSE
      gmul2(188) WHEN s_0_1 = to_unsigned(16#BD#, 8) ELSE
      gmul2(189) WHEN s_0_1 = to_unsigned(16#BE#, 8) ELSE
      gmul2(190) WHEN s_0_1 = to_unsigned(16#BF#, 8) ELSE
      gmul2(191) WHEN s_0_1 = to_unsigned(16#C0#, 8) ELSE
      gmul2(192) WHEN s_0_1 = to_unsigned(16#C1#, 8) ELSE
      gmul2(193) WHEN s_0_1 = to_unsigned(16#C2#, 8) ELSE
      gmul2(194) WHEN s_0_1 = to_unsigned(16#C3#, 8) ELSE
      gmul2(195) WHEN s_0_1 = to_unsigned(16#C4#, 8) ELSE
      gmul2(196) WHEN s_0_1 = to_unsigned(16#C5#, 8) ELSE
      gmul2(197) WHEN s_0_1 = to_unsigned(16#C6#, 8) ELSE
      gmul2(198) WHEN s_0_1 = to_unsigned(16#C7#, 8) ELSE
      gmul2(199) WHEN s_0_1 = to_unsigned(16#C8#, 8) ELSE
      gmul2(200) WHEN s_0_1 = to_unsigned(16#C9#, 8) ELSE
      gmul2(201) WHEN s_0_1 = to_unsigned(16#CA#, 8) ELSE
      gmul2(202) WHEN s_0_1 = to_unsigned(16#CB#, 8) ELSE
      gmul2(203) WHEN s_0_1 = to_unsigned(16#CC#, 8) ELSE
      gmul2(204) WHEN s_0_1 = to_unsigned(16#CD#, 8) ELSE
      gmul2(205) WHEN s_0_1 = to_unsigned(16#CE#, 8) ELSE
      gmul2(206) WHEN s_0_1 = to_unsigned(16#CF#, 8) ELSE
      gmul2(207) WHEN s_0_1 = to_unsigned(16#D0#, 8) ELSE
      gmul2(208) WHEN s_0_1 = to_unsigned(16#D1#, 8) ELSE
      gmul2(209) WHEN s_0_1 = to_unsigned(16#D2#, 8) ELSE
      gmul2(210) WHEN s_0_1 = to_unsigned(16#D3#, 8) ELSE
      gmul2(211) WHEN s_0_1 = to_unsigned(16#D4#, 8) ELSE
      gmul2(212) WHEN s_0_1 = to_unsigned(16#D5#, 8) ELSE
      gmul2(213) WHEN s_0_1 = to_unsigned(16#D6#, 8) ELSE
      gmul2(214) WHEN s_0_1 = to_unsigned(16#D7#, 8) ELSE
      gmul2(215) WHEN s_0_1 = to_unsigned(16#D8#, 8) ELSE
      gmul2(216) WHEN s_0_1 = to_unsigned(16#D9#, 8) ELSE
      gmul2(217) WHEN s_0_1 = to_unsigned(16#DA#, 8) ELSE
      gmul2(218) WHEN s_0_1 = to_unsigned(16#DB#, 8) ELSE
      gmul2(219) WHEN s_0_1 = to_unsigned(16#DC#, 8) ELSE
      gmul2(220) WHEN s_0_1 = to_unsigned(16#DD#, 8) ELSE
      gmul2(221) WHEN s_0_1 = to_unsigned(16#DE#, 8) ELSE
      gmul2(222) WHEN s_0_1 = to_unsigned(16#DF#, 8) ELSE
      gmul2(223) WHEN s_0_1 = to_unsigned(16#E0#, 8) ELSE
      gmul2(224) WHEN s_0_1 = to_unsigned(16#E1#, 8) ELSE
      gmul2(225) WHEN s_0_1 = to_unsigned(16#E2#, 8) ELSE
      gmul2(226) WHEN s_0_1 = to_unsigned(16#E3#, 8) ELSE
      gmul2(227) WHEN s_0_1 = to_unsigned(16#E4#, 8) ELSE
      gmul2(228) WHEN s_0_1 = to_unsigned(16#E5#, 8) ELSE
      gmul2(229) WHEN s_0_1 = to_unsigned(16#E6#, 8) ELSE
      gmul2(230) WHEN s_0_1 = to_unsigned(16#E7#, 8) ELSE
      gmul2(231) WHEN s_0_1 = to_unsigned(16#E8#, 8) ELSE
      gmul2(232) WHEN s_0_1 = to_unsigned(16#E9#, 8) ELSE
      gmul2(233) WHEN s_0_1 = to_unsigned(16#EA#, 8) ELSE
      gmul2(234) WHEN s_0_1 = to_unsigned(16#EB#, 8) ELSE
      gmul2(235) WHEN s_0_1 = to_unsigned(16#EC#, 8) ELSE
      gmul2(236) WHEN s_0_1 = to_unsigned(16#ED#, 8) ELSE
      gmul2(237) WHEN s_0_1 = to_unsigned(16#EE#, 8) ELSE
      gmul2(238) WHEN s_0_1 = to_unsigned(16#EF#, 8) ELSE
      gmul2(239) WHEN s_0_1 = to_unsigned(16#F0#, 8) ELSE
      gmul2(240) WHEN s_0_1 = to_unsigned(16#F1#, 8) ELSE
      gmul2(241) WHEN s_0_1 = to_unsigned(16#F2#, 8) ELSE
      gmul2(242) WHEN s_0_1 = to_unsigned(16#F3#, 8) ELSE
      gmul2(243) WHEN s_0_1 = to_unsigned(16#F4#, 8) ELSE
      gmul2(244) WHEN s_0_1 = to_unsigned(16#F5#, 8) ELSE
      gmul2(245) WHEN s_0_1 = to_unsigned(16#F6#, 8) ELSE
      gmul2(246) WHEN s_0_1 = to_unsigned(16#F7#, 8) ELSE
      gmul2(247) WHEN s_0_1 = to_unsigned(16#F8#, 8) ELSE
      gmul2(248) WHEN s_0_1 = to_unsigned(16#F9#, 8) ELSE
      gmul2(249) WHEN s_0_1 = to_unsigned(16#FA#, 8) ELSE
      gmul2(250) WHEN s_0_1 = to_unsigned(16#FB#, 8) ELSE
      gmul2(251) WHEN s_0_1 = to_unsigned(16#FC#, 8) ELSE
      gmul2(252) WHEN s_0_1 = to_unsigned(16#FD#, 8) ELSE
      gmul2(253) WHEN s_0_1 = to_unsigned(16#FE#, 8) ELSE
      gmul2(254) WHEN s_0_1 = to_unsigned(16#FF#, 8) ELSE
      gmul2(255);

  out0_189 <= out0_188 XOR out0_187;

  b1_3 <= out0_189 XOR s_2_1;

  out0_190 <= b1_3 XOR s_3_1;

  s_s_7(0) <= out0_190;
  s_s_7(1) <= s_s_1(1);
  s_s_7(2) <= s_s_1(2);
  s_s_7(3) <= s_s_1(3);
  s_s_7(4) <= s_s_1(4);
  s_s_7(5) <= s_s_1(5);
  s_s_7(6) <= s_s_1(6);
  s_s_7(7) <= s_s_1(7);
  s_s_7(8) <= s_s_1(8);
  s_s_7(9) <= s_s_1(9);
  s_s_7(10) <= s_s_1(10);
  s_s_7(11) <= s_s_1(11);
  s_s_7(12) <= s_s_1(12);
  s_s_7(13) <= s_s_1(13);
  s_s_7(14) <= s_s_1(14);
  s_s_7(15) <= s_s_1(15);

  s_s_8(0) <= s_s_7(0);
  s_s_8(1) <= out0_186;
  s_s_8(2) <= s_s_7(2);
  s_s_8(3) <= s_s_7(3);
  s_s_8(4) <= s_s_7(4);
  s_s_8(5) <= s_s_7(5);
  s_s_8(6) <= s_s_7(6);
  s_s_8(7) <= s_s_7(7);
  s_s_8(8) <= s_s_7(8);
  s_s_8(9) <= s_s_7(9);
  s_s_8(10) <= s_s_7(10);
  s_s_8(11) <= s_s_7(11);
  s_s_8(12) <= s_s_7(12);
  s_s_8(13) <= s_s_7(13);
  s_s_8(14) <= s_s_7(14);
  s_s_8(15) <= s_s_7(15);

  s_s_9(0) <= s_s_8(0);
  s_s_9(1) <= s_s_8(1);
  s_s_9(2) <= out0_182;
  s_s_9(3) <= s_s_8(3);
  s_s_9(4) <= s_s_8(4);
  s_s_9(5) <= s_s_8(5);
  s_s_9(6) <= s_s_8(6);
  s_s_9(7) <= s_s_8(7);
  s_s_9(8) <= s_s_8(8);
  s_s_9(9) <= s_s_8(9);
  s_s_9(10) <= s_s_8(10);
  s_s_9(11) <= s_s_8(11);
  s_s_9(12) <= s_s_8(12);
  s_s_9(13) <= s_s_8(13);
  s_s_9(14) <= s_s_8(14);
  s_s_9(15) <= s_s_8(15);

  s_s_6(0) <= s_s_9(0);
  s_s_6(1) <= s_s_9(1);
  s_s_6(2) <= s_s_9(2);
  s_s_6(3) <= out0_178;
  s_s_6(4) <= s_s_9(4);
  s_s_6(5) <= s_s_9(5);
  s_s_6(6) <= s_s_9(6);
  s_s_6(7) <= s_s_9(7);
  s_s_6(8) <= s_s_9(8);
  s_s_6(9) <= s_s_9(9);
  s_s_6(10) <= s_s_9(10);
  s_s_6(11) <= s_s_9(11);
  s_s_6(12) <= s_s_9(12);
  s_s_6(13) <= s_s_9(13);
  s_s_6(14) <= s_s_9(14);
  s_s_6(15) <= s_s_9(15);

  s_s_10(0) <= s_s_6(0);
  s_s_10(1) <= s_s_6(1);
  s_s_10(2) <= s_s_6(2);
  s_s_10(3) <= s_s_6(3);
  s_s_10(4) <= out0_174;
  s_s_10(5) <= s_s_6(5);
  s_s_10(6) <= s_s_6(6);
  s_s_10(7) <= s_s_6(7);
  s_s_10(8) <= s_s_6(8);
  s_s_10(9) <= s_s_6(9);
  s_s_10(10) <= s_s_6(10);
  s_s_10(11) <= s_s_6(11);
  s_s_10(12) <= s_s_6(12);
  s_s_10(13) <= s_s_6(13);
  s_s_10(14) <= s_s_6(14);
  s_s_10(15) <= s_s_6(15);

  s_s_11(0) <= s_s_10(0);
  s_s_11(1) <= s_s_10(1);
  s_s_11(2) <= s_s_10(2);
  s_s_11(3) <= s_s_10(3);
  s_s_11(4) <= s_s_10(4);
  s_s_11(5) <= out0_170;
  s_s_11(6) <= s_s_10(6);
  s_s_11(7) <= s_s_10(7);
  s_s_11(8) <= s_s_10(8);
  s_s_11(9) <= s_s_10(9);
  s_s_11(10) <= s_s_10(10);
  s_s_11(11) <= s_s_10(11);
  s_s_11(12) <= s_s_10(12);
  s_s_11(13) <= s_s_10(13);
  s_s_11(14) <= s_s_10(14);
  s_s_11(15) <= s_s_10(15);

  s_s_12(0) <= s_s_11(0);
  s_s_12(1) <= s_s_11(1);
  s_s_12(2) <= s_s_11(2);
  s_s_12(3) <= s_s_11(3);
  s_s_12(4) <= s_s_11(4);
  s_s_12(5) <= s_s_11(5);
  s_s_12(6) <= out0_166;
  s_s_12(7) <= s_s_11(7);
  s_s_12(8) <= s_s_11(8);
  s_s_12(9) <= s_s_11(9);
  s_s_12(10) <= s_s_11(10);
  s_s_12(11) <= s_s_11(11);
  s_s_12(12) <= s_s_11(12);
  s_s_12(13) <= s_s_11(13);
  s_s_12(14) <= s_s_11(14);
  s_s_12(15) <= s_s_11(15);

  s_s_5(0) <= s_s_12(0);
  s_s_5(1) <= s_s_12(1);
  s_s_5(2) <= s_s_12(2);
  s_s_5(3) <= s_s_12(3);
  s_s_5(4) <= s_s_12(4);
  s_s_5(5) <= s_s_12(5);
  s_s_5(6) <= s_s_12(6);
  s_s_5(7) <= out0_162;
  s_s_5(8) <= s_s_12(8);
  s_s_5(9) <= s_s_12(9);
  s_s_5(10) <= s_s_12(10);
  s_s_5(11) <= s_s_12(11);
  s_s_5(12) <= s_s_12(12);
  s_s_5(13) <= s_s_12(13);
  s_s_5(14) <= s_s_12(14);
  s_s_5(15) <= s_s_12(15);

  s_s_13(0) <= s_s_5(0);
  s_s_13(1) <= s_s_5(1);
  s_s_13(2) <= s_s_5(2);
  s_s_13(3) <= s_s_5(3);
  s_s_13(4) <= s_s_5(4);
  s_s_13(5) <= s_s_5(5);
  s_s_13(6) <= s_s_5(6);
  s_s_13(7) <= s_s_5(7);
  s_s_13(8) <= out0_158;
  s_s_13(9) <= s_s_5(9);
  s_s_13(10) <= s_s_5(10);
  s_s_13(11) <= s_s_5(11);
  s_s_13(12) <= s_s_5(12);
  s_s_13(13) <= s_s_5(13);
  s_s_13(14) <= s_s_5(14);
  s_s_13(15) <= s_s_5(15);

  s_s_14(0) <= s_s_13(0);
  s_s_14(1) <= s_s_13(1);
  s_s_14(2) <= s_s_13(2);
  s_s_14(3) <= s_s_13(3);
  s_s_14(4) <= s_s_13(4);
  s_s_14(5) <= s_s_13(5);
  s_s_14(6) <= s_s_13(6);
  s_s_14(7) <= s_s_13(7);
  s_s_14(8) <= s_s_13(8);
  s_s_14(9) <= out0_154;
  s_s_14(10) <= s_s_13(10);
  s_s_14(11) <= s_s_13(11);
  s_s_14(12) <= s_s_13(12);
  s_s_14(13) <= s_s_13(13);
  s_s_14(14) <= s_s_13(14);
  s_s_14(15) <= s_s_13(15);

  s_s_15(0) <= s_s_14(0);
  s_s_15(1) <= s_s_14(1);
  s_s_15(2) <= s_s_14(2);
  s_s_15(3) <= s_s_14(3);
  s_s_15(4) <= s_s_14(4);
  s_s_15(5) <= s_s_14(5);
  s_s_15(6) <= s_s_14(6);
  s_s_15(7) <= s_s_14(7);
  s_s_15(8) <= s_s_14(8);
  s_s_15(9) <= s_s_14(9);
  s_s_15(10) <= out0_150;
  s_s_15(11) <= s_s_14(11);
  s_s_15(12) <= s_s_14(12);
  s_s_15(13) <= s_s_14(13);
  s_s_15(14) <= s_s_14(14);
  s_s_15(15) <= s_s_14(15);

  s_s_4(0) <= s_s_15(0);
  s_s_4(1) <= s_s_15(1);
  s_s_4(2) <= s_s_15(2);
  s_s_4(3) <= s_s_15(3);
  s_s_4(4) <= s_s_15(4);
  s_s_4(5) <= s_s_15(5);
  s_s_4(6) <= s_s_15(6);
  s_s_4(7) <= s_s_15(7);
  s_s_4(8) <= s_s_15(8);
  s_s_4(9) <= s_s_15(9);
  s_s_4(10) <= s_s_15(10);
  s_s_4(11) <= out0_146;
  s_s_4(12) <= s_s_15(12);
  s_s_4(13) <= s_s_15(13);
  s_s_4(14) <= s_s_15(14);
  s_s_4(15) <= s_s_15(15);

  s_s_16(0) <= s_s_4(0);
  s_s_16(1) <= s_s_4(1);
  s_s_16(2) <= s_s_4(2);
  s_s_16(3) <= s_s_4(3);
  s_s_16(4) <= s_s_4(4);
  s_s_16(5) <= s_s_4(5);
  s_s_16(6) <= s_s_4(6);
  s_s_16(7) <= s_s_4(7);
  s_s_16(8) <= s_s_4(8);
  s_s_16(9) <= s_s_4(9);
  s_s_16(10) <= s_s_4(10);
  s_s_16(11) <= s_s_4(11);
  s_s_16(12) <= out0_142;
  s_s_16(13) <= s_s_4(13);
  s_s_16(14) <= s_s_4(14);
  s_s_16(15) <= s_s_4(15);

  s_s_17(0) <= s_s_16(0);
  s_s_17(1) <= s_s_16(1);
  s_s_17(2) <= s_s_16(2);
  s_s_17(3) <= s_s_16(3);
  s_s_17(4) <= s_s_16(4);
  s_s_17(5) <= s_s_16(5);
  s_s_17(6) <= s_s_16(6);
  s_s_17(7) <= s_s_16(7);
  s_s_17(8) <= s_s_16(8);
  s_s_17(9) <= s_s_16(9);
  s_s_17(10) <= s_s_16(10);
  s_s_17(11) <= s_s_16(11);
  s_s_17(12) <= s_s_16(12);
  s_s_17(13) <= out0_138;
  s_s_17(14) <= s_s_16(14);
  s_s_17(15) <= s_s_16(15);

  s_s_18(0) <= s_s_17(0);
  s_s_18(1) <= s_s_17(1);
  s_s_18(2) <= s_s_17(2);
  s_s_18(3) <= s_s_17(3);
  s_s_18(4) <= s_s_17(4);
  s_s_18(5) <= s_s_17(5);
  s_s_18(6) <= s_s_17(6);
  s_s_18(7) <= s_s_17(7);
  s_s_18(8) <= s_s_17(8);
  s_s_18(9) <= s_s_17(9);
  s_s_18(10) <= s_s_17(10);
  s_s_18(11) <= s_s_17(11);
  s_s_18(12) <= s_s_17(12);
  s_s_18(13) <= s_s_17(13);
  s_s_18(14) <= out0_134;
  s_s_18(15) <= s_s_17(15);

  s_s_19(0) <= s_s_18(0);
  s_s_19(1) <= s_s_18(1);
  s_s_19(2) <= s_s_18(2);
  s_s_19(3) <= s_s_18(3);
  s_s_19(4) <= s_s_18(4);
  s_s_19(5) <= s_s_18(5);
  s_s_19(6) <= s_s_18(6);
  s_s_19(7) <= s_s_18(7);
  s_s_19(8) <= s_s_18(8);
  s_s_19(9) <= s_s_18(9);
  s_s_19(10) <= s_s_18(10);
  s_s_19(11) <= s_s_18(11);
  s_s_19(12) <= s_s_18(12);
  s_s_19(13) <= s_s_18(13);
  s_s_19(14) <= s_s_18(14);
  s_s_19(15) <= out0_130;

  
  out0_191 <= s_s_1(0) WHEN ii_8 = to_unsigned(16#01#, 8) ELSE
      s_s_1(1) WHEN ii_8 = to_unsigned(16#02#, 8) ELSE
      s_s_1(2) WHEN ii_8 = to_unsigned(16#03#, 8) ELSE
      s_s_1(3) WHEN ii_8 = to_unsigned(16#04#, 8) ELSE
      s_s_1(4) WHEN ii_8 = to_unsigned(16#05#, 8) ELSE
      s_s_1(5) WHEN ii_8 = to_unsigned(16#06#, 8) ELSE
      s_s_1(6) WHEN ii_8 = to_unsigned(16#07#, 8) ELSE
      s_s_1(7) WHEN ii_8 = to_unsigned(16#08#, 8) ELSE
      s_s_1(8) WHEN ii_8 = to_unsigned(16#09#, 8) ELSE
      s_s_1(9) WHEN ii_8 = to_unsigned(16#0A#, 8) ELSE
      s_s_1(10) WHEN ii_8 = to_unsigned(16#0B#, 8) ELSE
      s_s_1(11) WHEN ii_8 = to_unsigned(16#0C#, 8) ELSE
      s_s_1(12) WHEN ii_8 = to_unsigned(16#0D#, 8) ELSE
      s_s_1(13) WHEN ii_8 = to_unsigned(16#0E#, 8) ELSE
      s_s_1(14) WHEN ii_8 = to_unsigned(16#0F#, 8) ELSE
      s_s_1(15);

  out0_192 <= out0_191 XOR out0_121;

  
  s_s_20(0) <= out0_192 WHEN ii_8 = to_unsigned(16#01#, 8) ELSE
      s_s_1(0);
  
  s_s_20(1) <= out0_192 WHEN ii_8 = to_unsigned(16#02#, 8) ELSE
      s_s_1(1);
  
  s_s_20(2) <= out0_192 WHEN ii_8 = to_unsigned(16#03#, 8) ELSE
      s_s_1(2);
  
  s_s_20(3) <= out0_192 WHEN ii_8 = to_unsigned(16#04#, 8) ELSE
      s_s_1(3);
  
  s_s_20(4) <= out0_192 WHEN ii_8 = to_unsigned(16#05#, 8) ELSE
      s_s_1(4);
  
  s_s_20(5) <= out0_192 WHEN ii_8 = to_unsigned(16#06#, 8) ELSE
      s_s_1(5);
  
  s_s_20(6) <= out0_192 WHEN ii_8 = to_unsigned(16#07#, 8) ELSE
      s_s_1(6);
  
  s_s_20(7) <= out0_192 WHEN ii_8 = to_unsigned(16#08#, 8) ELSE
      s_s_1(7);
  
  s_s_20(8) <= out0_192 WHEN ii_8 = to_unsigned(16#09#, 8) ELSE
      s_s_1(8);
  
  s_s_20(9) <= out0_192 WHEN ii_8 = to_unsigned(16#0A#, 8) ELSE
      s_s_1(9);
  
  s_s_20(10) <= out0_192 WHEN ii_8 = to_unsigned(16#0B#, 8) ELSE
      s_s_1(10);
  
  s_s_20(11) <= out0_192 WHEN ii_8 = to_unsigned(16#0C#, 8) ELSE
      s_s_1(11);
  
  s_s_20(12) <= out0_192 WHEN ii_8 = to_unsigned(16#0D#, 8) ELSE
      s_s_1(12);
  
  s_s_20(13) <= out0_192 WHEN ii_8 = to_unsigned(16#0E#, 8) ELSE
      s_s_1(13);
  
  s_s_20(14) <= out0_192 WHEN ii_8 = to_unsigned(16#0F#, 8) ELSE
      s_s_1(14);
  
  s_s_20(15) <= out0_192 WHEN ii_8 = to_unsigned(16#10#, 8) ELSE
      s_s_1(15);

  intdelay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        s_s_1(0) <= to_unsigned(16#00#, 8);
        s_s_1(1) <= to_unsigned(16#00#, 8);
        s_s_1(2) <= to_unsigned(16#00#, 8);
        s_s_1(3) <= to_unsigned(16#00#, 8);
        s_s_1(4) <= to_unsigned(16#00#, 8);
        s_s_1(5) <= to_unsigned(16#00#, 8);
        s_s_1(6) <= to_unsigned(16#00#, 8);
        s_s_1(7) <= to_unsigned(16#00#, 8);
        s_s_1(8) <= to_unsigned(16#00#, 8);
        s_s_1(9) <= to_unsigned(16#00#, 8);
        s_s_1(10) <= to_unsigned(16#00#, 8);
        s_s_1(11) <= to_unsigned(16#00#, 8);
        s_s_1(12) <= to_unsigned(16#00#, 8);
        s_s_1(13) <= to_unsigned(16#00#, 8);
        s_s_1(14) <= to_unsigned(16#00#, 8);
        s_s_1(15) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        s_s_1(0) <= s_s_21(0);
        s_s_1(1) <= s_s_21(1);
        s_s_1(2) <= s_s_21(2);
        s_s_1(3) <= s_s_21(3);
        s_s_1(4) <= s_s_21(4);
        s_s_1(5) <= s_s_21(5);
        s_s_1(6) <= s_s_21(6);
        s_s_1(7) <= s_s_21(7);
        s_s_1(8) <= s_s_21(8);
        s_s_1(9) <= s_s_21(9);
        s_s_1(10) <= s_s_21(10);
        s_s_1(11) <= s_s_21(11);
        s_s_1(12) <= s_s_21(12);
        s_s_1(13) <= s_s_21(13);
        s_s_1(14) <= s_s_21(14);
        s_s_1(15) <= s_s_21(15);
      END IF;
    END IF;
  END PROCESS intdelay3_process;


  
  out0_193(0) <= s_s_1(0) WHEN out0_10 = '0' ELSE
      s_s_1(0);
  
  out0_193(1) <= s_s_1(1) WHEN out0_10 = '0' ELSE
      s_s_1(1);
  
  out0_193(2) <= s_s_1(2) WHEN out0_10 = '0' ELSE
      s_s_1(2);
  
  out0_193(3) <= s_s_1(3) WHEN out0_10 = '0' ELSE
      s_s_1(3);
  
  out0_193(4) <= s_s_1(4) WHEN out0_10 = '0' ELSE
      s_s_1(4);
  
  out0_193(5) <= s_s_1(5) WHEN out0_10 = '0' ELSE
      s_s_1(5);
  
  out0_193(6) <= s_s_1(6) WHEN out0_10 = '0' ELSE
      s_s_1(6);
  
  out0_193(7) <= s_s_1(7) WHEN out0_10 = '0' ELSE
      s_s_1(7);
  
  out0_193(8) <= s_s_1(8) WHEN out0_10 = '0' ELSE
      s_s_1(8);
  
  out0_193(9) <= s_s_1(9) WHEN out0_10 = '0' ELSE
      s_s_1(9);
  
  out0_193(10) <= s_s_1(10) WHEN out0_10 = '0' ELSE
      s_s_1(10);
  
  out0_193(11) <= s_s_1(11) WHEN out0_10 = '0' ELSE
      s_s_1(11);
  
  out0_193(12) <= s_s_1(12) WHEN out0_10 = '0' ELSE
      s_s_1(12);
  
  out0_193(13) <= s_s_1(13) WHEN out0_10 = '0' ELSE
      s_s_1(13);
  
  out0_193(14) <= s_s_1(14) WHEN out0_10 = '0' ELSE
      s_s_1(14);
  
  out0_193(15) <= s_s_1(15) WHEN out0_10 = '0' ELSE
      s_s_1(15);

  
  out0_194(0) <= out0_193(0) WHEN out0_12 = '0' ELSE
      s_s_20(0);
  
  out0_194(1) <= out0_193(1) WHEN out0_12 = '0' ELSE
      s_s_20(1);
  
  out0_194(2) <= out0_193(2) WHEN out0_12 = '0' ELSE
      s_s_20(2);
  
  out0_194(3) <= out0_193(3) WHEN out0_12 = '0' ELSE
      s_s_20(3);
  
  out0_194(4) <= out0_193(4) WHEN out0_12 = '0' ELSE
      s_s_20(4);
  
  out0_194(5) <= out0_193(5) WHEN out0_12 = '0' ELSE
      s_s_20(5);
  
  out0_194(6) <= out0_193(6) WHEN out0_12 = '0' ELSE
      s_s_20(6);
  
  out0_194(7) <= out0_193(7) WHEN out0_12 = '0' ELSE
      s_s_20(7);
  
  out0_194(8) <= out0_193(8) WHEN out0_12 = '0' ELSE
      s_s_20(8);
  
  out0_194(9) <= out0_193(9) WHEN out0_12 = '0' ELSE
      s_s_20(9);
  
  out0_194(10) <= out0_193(10) WHEN out0_12 = '0' ELSE
      s_s_20(10);
  
  out0_194(11) <= out0_193(11) WHEN out0_12 = '0' ELSE
      s_s_20(11);
  
  out0_194(12) <= out0_193(12) WHEN out0_12 = '0' ELSE
      s_s_20(12);
  
  out0_194(13) <= out0_193(13) WHEN out0_12 = '0' ELSE
      s_s_20(13);
  
  out0_194(14) <= out0_193(14) WHEN out0_12 = '0' ELSE
      s_s_20(14);
  
  out0_194(15) <= out0_193(15) WHEN out0_12 = '0' ELSE
      s_s_20(15);

  
  out0_195(0) <= out0_194(0) WHEN out0_14 = '0' ELSE
      s_s_19(0);
  
  out0_195(1) <= out0_194(1) WHEN out0_14 = '0' ELSE
      s_s_19(1);
  
  out0_195(2) <= out0_194(2) WHEN out0_14 = '0' ELSE
      s_s_19(2);
  
  out0_195(3) <= out0_194(3) WHEN out0_14 = '0' ELSE
      s_s_19(3);
  
  out0_195(4) <= out0_194(4) WHEN out0_14 = '0' ELSE
      s_s_19(4);
  
  out0_195(5) <= out0_194(5) WHEN out0_14 = '0' ELSE
      s_s_19(5);
  
  out0_195(6) <= out0_194(6) WHEN out0_14 = '0' ELSE
      s_s_19(6);
  
  out0_195(7) <= out0_194(7) WHEN out0_14 = '0' ELSE
      s_s_19(7);
  
  out0_195(8) <= out0_194(8) WHEN out0_14 = '0' ELSE
      s_s_19(8);
  
  out0_195(9) <= out0_194(9) WHEN out0_14 = '0' ELSE
      s_s_19(9);
  
  out0_195(10) <= out0_194(10) WHEN out0_14 = '0' ELSE
      s_s_19(10);
  
  out0_195(11) <= out0_194(11) WHEN out0_14 = '0' ELSE
      s_s_19(11);
  
  out0_195(12) <= out0_194(12) WHEN out0_14 = '0' ELSE
      s_s_19(12);
  
  out0_195(13) <= out0_194(13) WHEN out0_14 = '0' ELSE
      s_s_19(13);
  
  out0_195(14) <= out0_194(14) WHEN out0_14 = '0' ELSE
      s_s_19(14);
  
  out0_195(15) <= out0_194(15) WHEN out0_14 = '0' ELSE
      s_s_19(15);

  
  out0_196(0) <= out0_195(0) WHEN out0_16 = '0' ELSE
      s_s_1(0);
  
  out0_196(1) <= out0_195(1) WHEN out0_16 = '0' ELSE
      s_s_1(1);
  
  out0_196(2) <= out0_195(2) WHEN out0_16 = '0' ELSE
      s_s_1(2);
  
  out0_196(3) <= out0_195(3) WHEN out0_16 = '0' ELSE
      s_s_1(3);
  
  out0_196(4) <= out0_195(4) WHEN out0_16 = '0' ELSE
      s_s_1(4);
  
  out0_196(5) <= out0_195(5) WHEN out0_16 = '0' ELSE
      s_s_1(5);
  
  out0_196(6) <= out0_195(6) WHEN out0_16 = '0' ELSE
      s_s_1(6);
  
  out0_196(7) <= out0_195(7) WHEN out0_16 = '0' ELSE
      s_s_1(7);
  
  out0_196(8) <= out0_195(8) WHEN out0_16 = '0' ELSE
      s_s_1(8);
  
  out0_196(9) <= out0_195(9) WHEN out0_16 = '0' ELSE
      s_s_1(9);
  
  out0_196(10) <= out0_195(10) WHEN out0_16 = '0' ELSE
      s_s_1(10);
  
  out0_196(11) <= out0_195(11) WHEN out0_16 = '0' ELSE
      s_s_1(11);
  
  out0_196(12) <= out0_195(12) WHEN out0_16 = '0' ELSE
      s_s_1(12);
  
  out0_196(13) <= out0_195(13) WHEN out0_16 = '0' ELSE
      s_s_1(13);
  
  out0_196(14) <= out0_195(14) WHEN out0_16 = '0' ELSE
      s_s_1(14);
  
  out0_196(15) <= out0_195(15) WHEN out0_16 = '0' ELSE
      s_s_1(15);

  
  out0_197(0) <= out0_196(0) WHEN out0_18 = '0' ELSE
      s_s_3(0);
  
  out0_197(1) <= out0_196(1) WHEN out0_18 = '0' ELSE
      s_s_3(1);
  
  out0_197(2) <= out0_196(2) WHEN out0_18 = '0' ELSE
      s_s_3(2);
  
  out0_197(3) <= out0_196(3) WHEN out0_18 = '0' ELSE
      s_s_3(3);
  
  out0_197(4) <= out0_196(4) WHEN out0_18 = '0' ELSE
      s_s_3(4);
  
  out0_197(5) <= out0_196(5) WHEN out0_18 = '0' ELSE
      s_s_3(5);
  
  out0_197(6) <= out0_196(6) WHEN out0_18 = '0' ELSE
      s_s_3(6);
  
  out0_197(7) <= out0_196(7) WHEN out0_18 = '0' ELSE
      s_s_3(7);
  
  out0_197(8) <= out0_196(8) WHEN out0_18 = '0' ELSE
      s_s_3(8);
  
  out0_197(9) <= out0_196(9) WHEN out0_18 = '0' ELSE
      s_s_3(9);
  
  out0_197(10) <= out0_196(10) WHEN out0_18 = '0' ELSE
      s_s_3(10);
  
  out0_197(11) <= out0_196(11) WHEN out0_18 = '0' ELSE
      s_s_3(11);
  
  out0_197(12) <= out0_196(12) WHEN out0_18 = '0' ELSE
      s_s_3(12);
  
  out0_197(13) <= out0_196(13) WHEN out0_18 = '0' ELSE
      s_s_3(13);
  
  out0_197(14) <= out0_196(14) WHEN out0_18 = '0' ELSE
      s_s_3(14);
  
  out0_197(15) <= out0_196(15) WHEN out0_18 = '0' ELSE
      s_s_3(15);

  
  out0_198(0) <= out0_197(0) WHEN out0_20 = '0' ELSE
      s_s_2(0);
  
  out0_198(1) <= out0_197(1) WHEN out0_20 = '0' ELSE
      s_s_2(1);
  
  out0_198(2) <= out0_197(2) WHEN out0_20 = '0' ELSE
      s_s_2(2);
  
  out0_198(3) <= out0_197(3) WHEN out0_20 = '0' ELSE
      s_s_2(3);
  
  out0_198(4) <= out0_197(4) WHEN out0_20 = '0' ELSE
      s_s_2(4);
  
  out0_198(5) <= out0_197(5) WHEN out0_20 = '0' ELSE
      s_s_2(5);
  
  out0_198(6) <= out0_197(6) WHEN out0_20 = '0' ELSE
      s_s_2(6);
  
  out0_198(7) <= out0_197(7) WHEN out0_20 = '0' ELSE
      s_s_2(7);
  
  out0_198(8) <= out0_197(8) WHEN out0_20 = '0' ELSE
      s_s_2(8);
  
  out0_198(9) <= out0_197(9) WHEN out0_20 = '0' ELSE
      s_s_2(9);
  
  out0_198(10) <= out0_197(10) WHEN out0_20 = '0' ELSE
      s_s_2(10);
  
  out0_198(11) <= out0_197(11) WHEN out0_20 = '0' ELSE
      s_s_2(11);
  
  out0_198(12) <= out0_197(12) WHEN out0_20 = '0' ELSE
      s_s_2(12);
  
  out0_198(13) <= out0_197(13) WHEN out0_20 = '0' ELSE
      s_s_2(13);
  
  out0_198(14) <= out0_197(14) WHEN out0_20 = '0' ELSE
      s_s_2(14);
  
  out0_198(15) <= out0_197(15) WHEN out0_20 = '0' ELSE
      s_s_2(15);

  
  out0_199(0) <= out0_198(0) WHEN out0_22 = '0' ELSE
      s_s_1(0);
  
  out0_199(1) <= out0_198(1) WHEN out0_22 = '0' ELSE
      s_s_1(1);
  
  out0_199(2) <= out0_198(2) WHEN out0_22 = '0' ELSE
      s_s_1(2);
  
  out0_199(3) <= out0_198(3) WHEN out0_22 = '0' ELSE
      s_s_1(3);
  
  out0_199(4) <= out0_198(4) WHEN out0_22 = '0' ELSE
      s_s_1(4);
  
  out0_199(5) <= out0_198(5) WHEN out0_22 = '0' ELSE
      s_s_1(5);
  
  out0_199(6) <= out0_198(6) WHEN out0_22 = '0' ELSE
      s_s_1(6);
  
  out0_199(7) <= out0_198(7) WHEN out0_22 = '0' ELSE
      s_s_1(7);
  
  out0_199(8) <= out0_198(8) WHEN out0_22 = '0' ELSE
      s_s_1(8);
  
  out0_199(9) <= out0_198(9) WHEN out0_22 = '0' ELSE
      s_s_1(9);
  
  out0_199(10) <= out0_198(10) WHEN out0_22 = '0' ELSE
      s_s_1(10);
  
  out0_199(11) <= out0_198(11) WHEN out0_22 = '0' ELSE
      s_s_1(11);
  
  out0_199(12) <= out0_198(12) WHEN out0_22 = '0' ELSE
      s_s_1(12);
  
  out0_199(13) <= out0_198(13) WHEN out0_22 = '0' ELSE
      s_s_1(13);
  
  out0_199(14) <= out0_198(14) WHEN out0_22 = '0' ELSE
      s_s_1(14);
  
  out0_199(15) <= out0_198(15) WHEN out0_22 = '0' ELSE
      s_s_1(15);

  
  s_s_21(0) <= out0_199(0) WHEN out0_24 = '0' ELSE
      s_s(0);
  
  s_s_21(1) <= out0_199(1) WHEN out0_24 = '0' ELSE
      s_s(1);
  
  s_s_21(2) <= out0_199(2) WHEN out0_24 = '0' ELSE
      s_s(2);
  
  s_s_21(3) <= out0_199(3) WHEN out0_24 = '0' ELSE
      s_s(3);
  
  s_s_21(4) <= out0_199(4) WHEN out0_24 = '0' ELSE
      s_s(4);
  
  s_s_21(5) <= out0_199(5) WHEN out0_24 = '0' ELSE
      s_s(5);
  
  s_s_21(6) <= out0_199(6) WHEN out0_24 = '0' ELSE
      s_s(6);
  
  s_s_21(7) <= out0_199(7) WHEN out0_24 = '0' ELSE
      s_s(7);
  
  s_s_21(8) <= out0_199(8) WHEN out0_24 = '0' ELSE
      s_s(8);
  
  s_s_21(9) <= out0_199(9) WHEN out0_24 = '0' ELSE
      s_s(9);
  
  s_s_21(10) <= out0_199(10) WHEN out0_24 = '0' ELSE
      s_s(10);
  
  s_s_21(11) <= out0_199(11) WHEN out0_24 = '0' ELSE
      s_s(11);
  
  s_s_21(12) <= out0_199(12) WHEN out0_24 = '0' ELSE
      s_s(12);
  
  s_s_21(13) <= out0_199(13) WHEN out0_24 = '0' ELSE
      s_s(13);
  
  s_s_21(14) <= out0_199(14) WHEN out0_24 = '0' ELSE
      s_s(14);
  
  s_s_21(15) <= out0_199(15) WHEN out0_24 = '0' ELSE
      s_s(15);

  Delay2_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay2_out1(0) <= to_unsigned(16#00#, 8);
        Delay2_out1(1) <= to_unsigned(16#00#, 8);
        Delay2_out1(2) <= to_unsigned(16#00#, 8);
        Delay2_out1(3) <= to_unsigned(16#00#, 8);
        Delay2_out1(4) <= to_unsigned(16#00#, 8);
        Delay2_out1(5) <= to_unsigned(16#00#, 8);
        Delay2_out1(6) <= to_unsigned(16#00#, 8);
        Delay2_out1(7) <= to_unsigned(16#00#, 8);
        Delay2_out1(8) <= to_unsigned(16#00#, 8);
        Delay2_out1(9) <= to_unsigned(16#00#, 8);
        Delay2_out1(10) <= to_unsigned(16#00#, 8);
        Delay2_out1(11) <= to_unsigned(16#00#, 8);
        Delay2_out1(12) <= to_unsigned(16#00#, 8);
        Delay2_out1(13) <= to_unsigned(16#00#, 8);
        Delay2_out1(14) <= to_unsigned(16#00#, 8);
        Delay2_out1(15) <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay2_out1(0) <= s_s_21(0);
        Delay2_out1(1) <= s_s_21(1);
        Delay2_out1(2) <= s_s_21(2);
        Delay2_out1(3) <= s_s_21(3);
        Delay2_out1(4) <= s_s_21(4);
        Delay2_out1(5) <= s_s_21(5);
        Delay2_out1(6) <= s_s_21(6);
        Delay2_out1(7) <= s_s_21(7);
        Delay2_out1(8) <= s_s_21(8);
        Delay2_out1(9) <= s_s_21(9);
        Delay2_out1(10) <= s_s_21(10);
        Delay2_out1(11) <= s_s_21(11);
        Delay2_out1(12) <= s_s_21(12);
        Delay2_out1(13) <= s_s_21(13);
        Delay2_out1(14) <= s_s_21(14);
        Delay2_out1(15) <= s_s_21(15);
      END IF;
    END IF;
  END PROCESS Delay2_process;


  outputgen: FOR kk IN 0 TO 15 GENERATE
    out_rsvd(kk) <= std_logic_vector(Delay2_out1(kk));
  END GENERATE;

  valid_1 <= to_unsigned(16#00#, 8);

  valid_2 <= to_unsigned(16#00#, 8);

  valid_3 <= to_unsigned(16#01#, 8);

  
  valid_4 <= valid_2 WHEN out0_40 = '0' ELSE
      valid_3;

  
  out0_200 <= valid_1 WHEN out0_10 = '0' ELSE
      valid_4;

  valid_5 <= to_unsigned(16#00#, 8);

  
  out0_201 <= out0_200 WHEN out0_12 = '0' ELSE
      valid_5;

  valid_6 <= to_unsigned(16#00#, 8);

  
  out0_202 <= out0_201 WHEN out0_14 = '0' ELSE
      valid_6;

  valid_7 <= to_unsigned(16#00#, 8);

  
  out0_203 <= out0_202 WHEN out0_16 = '0' ELSE
      valid_7;

  valid_8 <= to_unsigned(16#00#, 8);

  
  out0_204 <= out0_203 WHEN out0_18 = '0' ELSE
      valid_8;

  valid_9 <= to_unsigned(16#00#, 8);

  
  out0_205 <= out0_204 WHEN out0_20 = '0' ELSE
      valid_9;

  valid_10 <= to_unsigned(16#00#, 8);

  
  out0_206 <= out0_205 WHEN out0_22 = '0' ELSE
      valid_10;

  valid_11 <= to_unsigned(16#00#, 8);

  
  valid_12 <= out0_206 WHEN out0_24 = '0' ELSE
      valid_11;

  Delay3_process : PROCESS (clk)
  BEGIN
    IF clk'EVENT AND clk = '1' THEN
      IF reset_x = '1' THEN
        Delay3_out1 <= to_unsigned(16#00#, 8);
      ELSIF enb = '1' THEN
        Delay3_out1 <= valid_12;
      END IF;
    END IF;
  END PROCESS Delay3_process;


  valid <= std_logic_vector(Delay3_out1);

  sit_out <= std_logic_vector(sit_out_tmp);

  ce_out <= clk_enable;

END rtl;

